
module add_1506(
    input [1505:0] a_i_c,a_i_s,
    input [1505:0] b_i_c,b_i_s,
    output [1505:0] c_o,
    output [1505:0] s_o
);

wire [1505:0] p;
assign p = 1506'h2f49352b949f8f4812c7e263157738b15f6d37c9bfc0cd4914d536ce3542642d5cfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;

wire ha_c,ha_s,fa_c,fa_s;
wire [2:0] M;
wire [1505:0] c_t,s_t,c_t2,s_t2;
wire [1505:0] c_f,s_f;
wire [1505:0] corr_add;
wire [1506:0] c,s;

// FAs
    
fa fau_0_0(a_i_c[0],a_i_s[0],b_i_c[0],c_t[0],s_t[0]);
fa fau_0_1(a_i_c[1],a_i_s[1],b_i_c[1],c_t[1],s_t[1]);
fa fau_0_2(a_i_c[2],a_i_s[2],b_i_c[2],c_t[2],s_t[2]);
fa fau_0_3(a_i_c[3],a_i_s[3],b_i_c[3],c_t[3],s_t[3]);
fa fau_0_4(a_i_c[4],a_i_s[4],b_i_c[4],c_t[4],s_t[4]);
fa fau_0_5(a_i_c[5],a_i_s[5],b_i_c[5],c_t[5],s_t[5]);
fa fau_0_6(a_i_c[6],a_i_s[6],b_i_c[6],c_t[6],s_t[6]);
fa fau_0_7(a_i_c[7],a_i_s[7],b_i_c[7],c_t[7],s_t[7]);
fa fau_0_8(a_i_c[8],a_i_s[8],b_i_c[8],c_t[8],s_t[8]);
fa fau_0_9(a_i_c[9],a_i_s[9],b_i_c[9],c_t[9],s_t[9]);
fa fau_0_10(a_i_c[10],a_i_s[10],b_i_c[10],c_t[10],s_t[10]);
fa fau_0_11(a_i_c[11],a_i_s[11],b_i_c[11],c_t[11],s_t[11]);
fa fau_0_12(a_i_c[12],a_i_s[12],b_i_c[12],c_t[12],s_t[12]);
fa fau_0_13(a_i_c[13],a_i_s[13],b_i_c[13],c_t[13],s_t[13]);
fa fau_0_14(a_i_c[14],a_i_s[14],b_i_c[14],c_t[14],s_t[14]);
fa fau_0_15(a_i_c[15],a_i_s[15],b_i_c[15],c_t[15],s_t[15]);
fa fau_0_16(a_i_c[16],a_i_s[16],b_i_c[16],c_t[16],s_t[16]);
fa fau_0_17(a_i_c[17],a_i_s[17],b_i_c[17],c_t[17],s_t[17]);
fa fau_0_18(a_i_c[18],a_i_s[18],b_i_c[18],c_t[18],s_t[18]);
fa fau_0_19(a_i_c[19],a_i_s[19],b_i_c[19],c_t[19],s_t[19]);
fa fau_0_20(a_i_c[20],a_i_s[20],b_i_c[20],c_t[20],s_t[20]);
fa fau_0_21(a_i_c[21],a_i_s[21],b_i_c[21],c_t[21],s_t[21]);
fa fau_0_22(a_i_c[22],a_i_s[22],b_i_c[22],c_t[22],s_t[22]);
fa fau_0_23(a_i_c[23],a_i_s[23],b_i_c[23],c_t[23],s_t[23]);
fa fau_0_24(a_i_c[24],a_i_s[24],b_i_c[24],c_t[24],s_t[24]);
fa fau_0_25(a_i_c[25],a_i_s[25],b_i_c[25],c_t[25],s_t[25]);
fa fau_0_26(a_i_c[26],a_i_s[26],b_i_c[26],c_t[26],s_t[26]);
fa fau_0_27(a_i_c[27],a_i_s[27],b_i_c[27],c_t[27],s_t[27]);
fa fau_0_28(a_i_c[28],a_i_s[28],b_i_c[28],c_t[28],s_t[28]);
fa fau_0_29(a_i_c[29],a_i_s[29],b_i_c[29],c_t[29],s_t[29]);
fa fau_0_30(a_i_c[30],a_i_s[30],b_i_c[30],c_t[30],s_t[30]);
fa fau_0_31(a_i_c[31],a_i_s[31],b_i_c[31],c_t[31],s_t[31]);
fa fau_0_32(a_i_c[32],a_i_s[32],b_i_c[32],c_t[32],s_t[32]);
fa fau_0_33(a_i_c[33],a_i_s[33],b_i_c[33],c_t[33],s_t[33]);
fa fau_0_34(a_i_c[34],a_i_s[34],b_i_c[34],c_t[34],s_t[34]);
fa fau_0_35(a_i_c[35],a_i_s[35],b_i_c[35],c_t[35],s_t[35]);
fa fau_0_36(a_i_c[36],a_i_s[36],b_i_c[36],c_t[36],s_t[36]);
fa fau_0_37(a_i_c[37],a_i_s[37],b_i_c[37],c_t[37],s_t[37]);
fa fau_0_38(a_i_c[38],a_i_s[38],b_i_c[38],c_t[38],s_t[38]);
fa fau_0_39(a_i_c[39],a_i_s[39],b_i_c[39],c_t[39],s_t[39]);
fa fau_0_40(a_i_c[40],a_i_s[40],b_i_c[40],c_t[40],s_t[40]);
fa fau_0_41(a_i_c[41],a_i_s[41],b_i_c[41],c_t[41],s_t[41]);
fa fau_0_42(a_i_c[42],a_i_s[42],b_i_c[42],c_t[42],s_t[42]);
fa fau_0_43(a_i_c[43],a_i_s[43],b_i_c[43],c_t[43],s_t[43]);
fa fau_0_44(a_i_c[44],a_i_s[44],b_i_c[44],c_t[44],s_t[44]);
fa fau_0_45(a_i_c[45],a_i_s[45],b_i_c[45],c_t[45],s_t[45]);
fa fau_0_46(a_i_c[46],a_i_s[46],b_i_c[46],c_t[46],s_t[46]);
fa fau_0_47(a_i_c[47],a_i_s[47],b_i_c[47],c_t[47],s_t[47]);
fa fau_0_48(a_i_c[48],a_i_s[48],b_i_c[48],c_t[48],s_t[48]);
fa fau_0_49(a_i_c[49],a_i_s[49],b_i_c[49],c_t[49],s_t[49]);
fa fau_0_50(a_i_c[50],a_i_s[50],b_i_c[50],c_t[50],s_t[50]);
fa fau_0_51(a_i_c[51],a_i_s[51],b_i_c[51],c_t[51],s_t[51]);
fa fau_0_52(a_i_c[52],a_i_s[52],b_i_c[52],c_t[52],s_t[52]);
fa fau_0_53(a_i_c[53],a_i_s[53],b_i_c[53],c_t[53],s_t[53]);
fa fau_0_54(a_i_c[54],a_i_s[54],b_i_c[54],c_t[54],s_t[54]);
fa fau_0_55(a_i_c[55],a_i_s[55],b_i_c[55],c_t[55],s_t[55]);
fa fau_0_56(a_i_c[56],a_i_s[56],b_i_c[56],c_t[56],s_t[56]);
fa fau_0_57(a_i_c[57],a_i_s[57],b_i_c[57],c_t[57],s_t[57]);
fa fau_0_58(a_i_c[58],a_i_s[58],b_i_c[58],c_t[58],s_t[58]);
fa fau_0_59(a_i_c[59],a_i_s[59],b_i_c[59],c_t[59],s_t[59]);
fa fau_0_60(a_i_c[60],a_i_s[60],b_i_c[60],c_t[60],s_t[60]);
fa fau_0_61(a_i_c[61],a_i_s[61],b_i_c[61],c_t[61],s_t[61]);
fa fau_0_62(a_i_c[62],a_i_s[62],b_i_c[62],c_t[62],s_t[62]);
fa fau_0_63(a_i_c[63],a_i_s[63],b_i_c[63],c_t[63],s_t[63]);
fa fau_0_64(a_i_c[64],a_i_s[64],b_i_c[64],c_t[64],s_t[64]);
fa fau_0_65(a_i_c[65],a_i_s[65],b_i_c[65],c_t[65],s_t[65]);
fa fau_0_66(a_i_c[66],a_i_s[66],b_i_c[66],c_t[66],s_t[66]);
fa fau_0_67(a_i_c[67],a_i_s[67],b_i_c[67],c_t[67],s_t[67]);
fa fau_0_68(a_i_c[68],a_i_s[68],b_i_c[68],c_t[68],s_t[68]);
fa fau_0_69(a_i_c[69],a_i_s[69],b_i_c[69],c_t[69],s_t[69]);
fa fau_0_70(a_i_c[70],a_i_s[70],b_i_c[70],c_t[70],s_t[70]);
fa fau_0_71(a_i_c[71],a_i_s[71],b_i_c[71],c_t[71],s_t[71]);
fa fau_0_72(a_i_c[72],a_i_s[72],b_i_c[72],c_t[72],s_t[72]);
fa fau_0_73(a_i_c[73],a_i_s[73],b_i_c[73],c_t[73],s_t[73]);
fa fau_0_74(a_i_c[74],a_i_s[74],b_i_c[74],c_t[74],s_t[74]);
fa fau_0_75(a_i_c[75],a_i_s[75],b_i_c[75],c_t[75],s_t[75]);
fa fau_0_76(a_i_c[76],a_i_s[76],b_i_c[76],c_t[76],s_t[76]);
fa fau_0_77(a_i_c[77],a_i_s[77],b_i_c[77],c_t[77],s_t[77]);
fa fau_0_78(a_i_c[78],a_i_s[78],b_i_c[78],c_t[78],s_t[78]);
fa fau_0_79(a_i_c[79],a_i_s[79],b_i_c[79],c_t[79],s_t[79]);
fa fau_0_80(a_i_c[80],a_i_s[80],b_i_c[80],c_t[80],s_t[80]);
fa fau_0_81(a_i_c[81],a_i_s[81],b_i_c[81],c_t[81],s_t[81]);
fa fau_0_82(a_i_c[82],a_i_s[82],b_i_c[82],c_t[82],s_t[82]);
fa fau_0_83(a_i_c[83],a_i_s[83],b_i_c[83],c_t[83],s_t[83]);
fa fau_0_84(a_i_c[84],a_i_s[84],b_i_c[84],c_t[84],s_t[84]);
fa fau_0_85(a_i_c[85],a_i_s[85],b_i_c[85],c_t[85],s_t[85]);
fa fau_0_86(a_i_c[86],a_i_s[86],b_i_c[86],c_t[86],s_t[86]);
fa fau_0_87(a_i_c[87],a_i_s[87],b_i_c[87],c_t[87],s_t[87]);
fa fau_0_88(a_i_c[88],a_i_s[88],b_i_c[88],c_t[88],s_t[88]);
fa fau_0_89(a_i_c[89],a_i_s[89],b_i_c[89],c_t[89],s_t[89]);
fa fau_0_90(a_i_c[90],a_i_s[90],b_i_c[90],c_t[90],s_t[90]);
fa fau_0_91(a_i_c[91],a_i_s[91],b_i_c[91],c_t[91],s_t[91]);
fa fau_0_92(a_i_c[92],a_i_s[92],b_i_c[92],c_t[92],s_t[92]);
fa fau_0_93(a_i_c[93],a_i_s[93],b_i_c[93],c_t[93],s_t[93]);
fa fau_0_94(a_i_c[94],a_i_s[94],b_i_c[94],c_t[94],s_t[94]);
fa fau_0_95(a_i_c[95],a_i_s[95],b_i_c[95],c_t[95],s_t[95]);
fa fau_0_96(a_i_c[96],a_i_s[96],b_i_c[96],c_t[96],s_t[96]);
fa fau_0_97(a_i_c[97],a_i_s[97],b_i_c[97],c_t[97],s_t[97]);
fa fau_0_98(a_i_c[98],a_i_s[98],b_i_c[98],c_t[98],s_t[98]);
fa fau_0_99(a_i_c[99],a_i_s[99],b_i_c[99],c_t[99],s_t[99]);
fa fau_0_100(a_i_c[100],a_i_s[100],b_i_c[100],c_t[100],s_t[100]);
fa fau_0_101(a_i_c[101],a_i_s[101],b_i_c[101],c_t[101],s_t[101]);
fa fau_0_102(a_i_c[102],a_i_s[102],b_i_c[102],c_t[102],s_t[102]);
fa fau_0_103(a_i_c[103],a_i_s[103],b_i_c[103],c_t[103],s_t[103]);
fa fau_0_104(a_i_c[104],a_i_s[104],b_i_c[104],c_t[104],s_t[104]);
fa fau_0_105(a_i_c[105],a_i_s[105],b_i_c[105],c_t[105],s_t[105]);
fa fau_0_106(a_i_c[106],a_i_s[106],b_i_c[106],c_t[106],s_t[106]);
fa fau_0_107(a_i_c[107],a_i_s[107],b_i_c[107],c_t[107],s_t[107]);
fa fau_0_108(a_i_c[108],a_i_s[108],b_i_c[108],c_t[108],s_t[108]);
fa fau_0_109(a_i_c[109],a_i_s[109],b_i_c[109],c_t[109],s_t[109]);
fa fau_0_110(a_i_c[110],a_i_s[110],b_i_c[110],c_t[110],s_t[110]);
fa fau_0_111(a_i_c[111],a_i_s[111],b_i_c[111],c_t[111],s_t[111]);
fa fau_0_112(a_i_c[112],a_i_s[112],b_i_c[112],c_t[112],s_t[112]);
fa fau_0_113(a_i_c[113],a_i_s[113],b_i_c[113],c_t[113],s_t[113]);
fa fau_0_114(a_i_c[114],a_i_s[114],b_i_c[114],c_t[114],s_t[114]);
fa fau_0_115(a_i_c[115],a_i_s[115],b_i_c[115],c_t[115],s_t[115]);
fa fau_0_116(a_i_c[116],a_i_s[116],b_i_c[116],c_t[116],s_t[116]);
fa fau_0_117(a_i_c[117],a_i_s[117],b_i_c[117],c_t[117],s_t[117]);
fa fau_0_118(a_i_c[118],a_i_s[118],b_i_c[118],c_t[118],s_t[118]);
fa fau_0_119(a_i_c[119],a_i_s[119],b_i_c[119],c_t[119],s_t[119]);
fa fau_0_120(a_i_c[120],a_i_s[120],b_i_c[120],c_t[120],s_t[120]);
fa fau_0_121(a_i_c[121],a_i_s[121],b_i_c[121],c_t[121],s_t[121]);
fa fau_0_122(a_i_c[122],a_i_s[122],b_i_c[122],c_t[122],s_t[122]);
fa fau_0_123(a_i_c[123],a_i_s[123],b_i_c[123],c_t[123],s_t[123]);
fa fau_0_124(a_i_c[124],a_i_s[124],b_i_c[124],c_t[124],s_t[124]);
fa fau_0_125(a_i_c[125],a_i_s[125],b_i_c[125],c_t[125],s_t[125]);
fa fau_0_126(a_i_c[126],a_i_s[126],b_i_c[126],c_t[126],s_t[126]);
fa fau_0_127(a_i_c[127],a_i_s[127],b_i_c[127],c_t[127],s_t[127]);
fa fau_0_128(a_i_c[128],a_i_s[128],b_i_c[128],c_t[128],s_t[128]);
fa fau_0_129(a_i_c[129],a_i_s[129],b_i_c[129],c_t[129],s_t[129]);
fa fau_0_130(a_i_c[130],a_i_s[130],b_i_c[130],c_t[130],s_t[130]);
fa fau_0_131(a_i_c[131],a_i_s[131],b_i_c[131],c_t[131],s_t[131]);
fa fau_0_132(a_i_c[132],a_i_s[132],b_i_c[132],c_t[132],s_t[132]);
fa fau_0_133(a_i_c[133],a_i_s[133],b_i_c[133],c_t[133],s_t[133]);
fa fau_0_134(a_i_c[134],a_i_s[134],b_i_c[134],c_t[134],s_t[134]);
fa fau_0_135(a_i_c[135],a_i_s[135],b_i_c[135],c_t[135],s_t[135]);
fa fau_0_136(a_i_c[136],a_i_s[136],b_i_c[136],c_t[136],s_t[136]);
fa fau_0_137(a_i_c[137],a_i_s[137],b_i_c[137],c_t[137],s_t[137]);
fa fau_0_138(a_i_c[138],a_i_s[138],b_i_c[138],c_t[138],s_t[138]);
fa fau_0_139(a_i_c[139],a_i_s[139],b_i_c[139],c_t[139],s_t[139]);
fa fau_0_140(a_i_c[140],a_i_s[140],b_i_c[140],c_t[140],s_t[140]);
fa fau_0_141(a_i_c[141],a_i_s[141],b_i_c[141],c_t[141],s_t[141]);
fa fau_0_142(a_i_c[142],a_i_s[142],b_i_c[142],c_t[142],s_t[142]);
fa fau_0_143(a_i_c[143],a_i_s[143],b_i_c[143],c_t[143],s_t[143]);
fa fau_0_144(a_i_c[144],a_i_s[144],b_i_c[144],c_t[144],s_t[144]);
fa fau_0_145(a_i_c[145],a_i_s[145],b_i_c[145],c_t[145],s_t[145]);
fa fau_0_146(a_i_c[146],a_i_s[146],b_i_c[146],c_t[146],s_t[146]);
fa fau_0_147(a_i_c[147],a_i_s[147],b_i_c[147],c_t[147],s_t[147]);
fa fau_0_148(a_i_c[148],a_i_s[148],b_i_c[148],c_t[148],s_t[148]);
fa fau_0_149(a_i_c[149],a_i_s[149],b_i_c[149],c_t[149],s_t[149]);
fa fau_0_150(a_i_c[150],a_i_s[150],b_i_c[150],c_t[150],s_t[150]);
fa fau_0_151(a_i_c[151],a_i_s[151],b_i_c[151],c_t[151],s_t[151]);
fa fau_0_152(a_i_c[152],a_i_s[152],b_i_c[152],c_t[152],s_t[152]);
fa fau_0_153(a_i_c[153],a_i_s[153],b_i_c[153],c_t[153],s_t[153]);
fa fau_0_154(a_i_c[154],a_i_s[154],b_i_c[154],c_t[154],s_t[154]);
fa fau_0_155(a_i_c[155],a_i_s[155],b_i_c[155],c_t[155],s_t[155]);
fa fau_0_156(a_i_c[156],a_i_s[156],b_i_c[156],c_t[156],s_t[156]);
fa fau_0_157(a_i_c[157],a_i_s[157],b_i_c[157],c_t[157],s_t[157]);
fa fau_0_158(a_i_c[158],a_i_s[158],b_i_c[158],c_t[158],s_t[158]);
fa fau_0_159(a_i_c[159],a_i_s[159],b_i_c[159],c_t[159],s_t[159]);
fa fau_0_160(a_i_c[160],a_i_s[160],b_i_c[160],c_t[160],s_t[160]);
fa fau_0_161(a_i_c[161],a_i_s[161],b_i_c[161],c_t[161],s_t[161]);
fa fau_0_162(a_i_c[162],a_i_s[162],b_i_c[162],c_t[162],s_t[162]);
fa fau_0_163(a_i_c[163],a_i_s[163],b_i_c[163],c_t[163],s_t[163]);
fa fau_0_164(a_i_c[164],a_i_s[164],b_i_c[164],c_t[164],s_t[164]);
fa fau_0_165(a_i_c[165],a_i_s[165],b_i_c[165],c_t[165],s_t[165]);
fa fau_0_166(a_i_c[166],a_i_s[166],b_i_c[166],c_t[166],s_t[166]);
fa fau_0_167(a_i_c[167],a_i_s[167],b_i_c[167],c_t[167],s_t[167]);
fa fau_0_168(a_i_c[168],a_i_s[168],b_i_c[168],c_t[168],s_t[168]);
fa fau_0_169(a_i_c[169],a_i_s[169],b_i_c[169],c_t[169],s_t[169]);
fa fau_0_170(a_i_c[170],a_i_s[170],b_i_c[170],c_t[170],s_t[170]);
fa fau_0_171(a_i_c[171],a_i_s[171],b_i_c[171],c_t[171],s_t[171]);
fa fau_0_172(a_i_c[172],a_i_s[172],b_i_c[172],c_t[172],s_t[172]);
fa fau_0_173(a_i_c[173],a_i_s[173],b_i_c[173],c_t[173],s_t[173]);
fa fau_0_174(a_i_c[174],a_i_s[174],b_i_c[174],c_t[174],s_t[174]);
fa fau_0_175(a_i_c[175],a_i_s[175],b_i_c[175],c_t[175],s_t[175]);
fa fau_0_176(a_i_c[176],a_i_s[176],b_i_c[176],c_t[176],s_t[176]);
fa fau_0_177(a_i_c[177],a_i_s[177],b_i_c[177],c_t[177],s_t[177]);
fa fau_0_178(a_i_c[178],a_i_s[178],b_i_c[178],c_t[178],s_t[178]);
fa fau_0_179(a_i_c[179],a_i_s[179],b_i_c[179],c_t[179],s_t[179]);
fa fau_0_180(a_i_c[180],a_i_s[180],b_i_c[180],c_t[180],s_t[180]);
fa fau_0_181(a_i_c[181],a_i_s[181],b_i_c[181],c_t[181],s_t[181]);
fa fau_0_182(a_i_c[182],a_i_s[182],b_i_c[182],c_t[182],s_t[182]);
fa fau_0_183(a_i_c[183],a_i_s[183],b_i_c[183],c_t[183],s_t[183]);
fa fau_0_184(a_i_c[184],a_i_s[184],b_i_c[184],c_t[184],s_t[184]);
fa fau_0_185(a_i_c[185],a_i_s[185],b_i_c[185],c_t[185],s_t[185]);
fa fau_0_186(a_i_c[186],a_i_s[186],b_i_c[186],c_t[186],s_t[186]);
fa fau_0_187(a_i_c[187],a_i_s[187],b_i_c[187],c_t[187],s_t[187]);
fa fau_0_188(a_i_c[188],a_i_s[188],b_i_c[188],c_t[188],s_t[188]);
fa fau_0_189(a_i_c[189],a_i_s[189],b_i_c[189],c_t[189],s_t[189]);
fa fau_0_190(a_i_c[190],a_i_s[190],b_i_c[190],c_t[190],s_t[190]);
fa fau_0_191(a_i_c[191],a_i_s[191],b_i_c[191],c_t[191],s_t[191]);
fa fau_0_192(a_i_c[192],a_i_s[192],b_i_c[192],c_t[192],s_t[192]);
fa fau_0_193(a_i_c[193],a_i_s[193],b_i_c[193],c_t[193],s_t[193]);
fa fau_0_194(a_i_c[194],a_i_s[194],b_i_c[194],c_t[194],s_t[194]);
fa fau_0_195(a_i_c[195],a_i_s[195],b_i_c[195],c_t[195],s_t[195]);
fa fau_0_196(a_i_c[196],a_i_s[196],b_i_c[196],c_t[196],s_t[196]);
fa fau_0_197(a_i_c[197],a_i_s[197],b_i_c[197],c_t[197],s_t[197]);
fa fau_0_198(a_i_c[198],a_i_s[198],b_i_c[198],c_t[198],s_t[198]);
fa fau_0_199(a_i_c[199],a_i_s[199],b_i_c[199],c_t[199],s_t[199]);
fa fau_0_200(a_i_c[200],a_i_s[200],b_i_c[200],c_t[200],s_t[200]);
fa fau_0_201(a_i_c[201],a_i_s[201],b_i_c[201],c_t[201],s_t[201]);
fa fau_0_202(a_i_c[202],a_i_s[202],b_i_c[202],c_t[202],s_t[202]);
fa fau_0_203(a_i_c[203],a_i_s[203],b_i_c[203],c_t[203],s_t[203]);
fa fau_0_204(a_i_c[204],a_i_s[204],b_i_c[204],c_t[204],s_t[204]);
fa fau_0_205(a_i_c[205],a_i_s[205],b_i_c[205],c_t[205],s_t[205]);
fa fau_0_206(a_i_c[206],a_i_s[206],b_i_c[206],c_t[206],s_t[206]);
fa fau_0_207(a_i_c[207],a_i_s[207],b_i_c[207],c_t[207],s_t[207]);
fa fau_0_208(a_i_c[208],a_i_s[208],b_i_c[208],c_t[208],s_t[208]);
fa fau_0_209(a_i_c[209],a_i_s[209],b_i_c[209],c_t[209],s_t[209]);
fa fau_0_210(a_i_c[210],a_i_s[210],b_i_c[210],c_t[210],s_t[210]);
fa fau_0_211(a_i_c[211],a_i_s[211],b_i_c[211],c_t[211],s_t[211]);
fa fau_0_212(a_i_c[212],a_i_s[212],b_i_c[212],c_t[212],s_t[212]);
fa fau_0_213(a_i_c[213],a_i_s[213],b_i_c[213],c_t[213],s_t[213]);
fa fau_0_214(a_i_c[214],a_i_s[214],b_i_c[214],c_t[214],s_t[214]);
fa fau_0_215(a_i_c[215],a_i_s[215],b_i_c[215],c_t[215],s_t[215]);
fa fau_0_216(a_i_c[216],a_i_s[216],b_i_c[216],c_t[216],s_t[216]);
fa fau_0_217(a_i_c[217],a_i_s[217],b_i_c[217],c_t[217],s_t[217]);
fa fau_0_218(a_i_c[218],a_i_s[218],b_i_c[218],c_t[218],s_t[218]);
fa fau_0_219(a_i_c[219],a_i_s[219],b_i_c[219],c_t[219],s_t[219]);
fa fau_0_220(a_i_c[220],a_i_s[220],b_i_c[220],c_t[220],s_t[220]);
fa fau_0_221(a_i_c[221],a_i_s[221],b_i_c[221],c_t[221],s_t[221]);
fa fau_0_222(a_i_c[222],a_i_s[222],b_i_c[222],c_t[222],s_t[222]);
fa fau_0_223(a_i_c[223],a_i_s[223],b_i_c[223],c_t[223],s_t[223]);
fa fau_0_224(a_i_c[224],a_i_s[224],b_i_c[224],c_t[224],s_t[224]);
fa fau_0_225(a_i_c[225],a_i_s[225],b_i_c[225],c_t[225],s_t[225]);
fa fau_0_226(a_i_c[226],a_i_s[226],b_i_c[226],c_t[226],s_t[226]);
fa fau_0_227(a_i_c[227],a_i_s[227],b_i_c[227],c_t[227],s_t[227]);
fa fau_0_228(a_i_c[228],a_i_s[228],b_i_c[228],c_t[228],s_t[228]);
fa fau_0_229(a_i_c[229],a_i_s[229],b_i_c[229],c_t[229],s_t[229]);
fa fau_0_230(a_i_c[230],a_i_s[230],b_i_c[230],c_t[230],s_t[230]);
fa fau_0_231(a_i_c[231],a_i_s[231],b_i_c[231],c_t[231],s_t[231]);
fa fau_0_232(a_i_c[232],a_i_s[232],b_i_c[232],c_t[232],s_t[232]);
fa fau_0_233(a_i_c[233],a_i_s[233],b_i_c[233],c_t[233],s_t[233]);
fa fau_0_234(a_i_c[234],a_i_s[234],b_i_c[234],c_t[234],s_t[234]);
fa fau_0_235(a_i_c[235],a_i_s[235],b_i_c[235],c_t[235],s_t[235]);
fa fau_0_236(a_i_c[236],a_i_s[236],b_i_c[236],c_t[236],s_t[236]);
fa fau_0_237(a_i_c[237],a_i_s[237],b_i_c[237],c_t[237],s_t[237]);
fa fau_0_238(a_i_c[238],a_i_s[238],b_i_c[238],c_t[238],s_t[238]);
fa fau_0_239(a_i_c[239],a_i_s[239],b_i_c[239],c_t[239],s_t[239]);
fa fau_0_240(a_i_c[240],a_i_s[240],b_i_c[240],c_t[240],s_t[240]);
fa fau_0_241(a_i_c[241],a_i_s[241],b_i_c[241],c_t[241],s_t[241]);
fa fau_0_242(a_i_c[242],a_i_s[242],b_i_c[242],c_t[242],s_t[242]);
fa fau_0_243(a_i_c[243],a_i_s[243],b_i_c[243],c_t[243],s_t[243]);
fa fau_0_244(a_i_c[244],a_i_s[244],b_i_c[244],c_t[244],s_t[244]);
fa fau_0_245(a_i_c[245],a_i_s[245],b_i_c[245],c_t[245],s_t[245]);
fa fau_0_246(a_i_c[246],a_i_s[246],b_i_c[246],c_t[246],s_t[246]);
fa fau_0_247(a_i_c[247],a_i_s[247],b_i_c[247],c_t[247],s_t[247]);
fa fau_0_248(a_i_c[248],a_i_s[248],b_i_c[248],c_t[248],s_t[248]);
fa fau_0_249(a_i_c[249],a_i_s[249],b_i_c[249],c_t[249],s_t[249]);
fa fau_0_250(a_i_c[250],a_i_s[250],b_i_c[250],c_t[250],s_t[250]);
fa fau_0_251(a_i_c[251],a_i_s[251],b_i_c[251],c_t[251],s_t[251]);
fa fau_0_252(a_i_c[252],a_i_s[252],b_i_c[252],c_t[252],s_t[252]);
fa fau_0_253(a_i_c[253],a_i_s[253],b_i_c[253],c_t[253],s_t[253]);
fa fau_0_254(a_i_c[254],a_i_s[254],b_i_c[254],c_t[254],s_t[254]);
fa fau_0_255(a_i_c[255],a_i_s[255],b_i_c[255],c_t[255],s_t[255]);
fa fau_0_256(a_i_c[256],a_i_s[256],b_i_c[256],c_t[256],s_t[256]);
fa fau_0_257(a_i_c[257],a_i_s[257],b_i_c[257],c_t[257],s_t[257]);
fa fau_0_258(a_i_c[258],a_i_s[258],b_i_c[258],c_t[258],s_t[258]);
fa fau_0_259(a_i_c[259],a_i_s[259],b_i_c[259],c_t[259],s_t[259]);
fa fau_0_260(a_i_c[260],a_i_s[260],b_i_c[260],c_t[260],s_t[260]);
fa fau_0_261(a_i_c[261],a_i_s[261],b_i_c[261],c_t[261],s_t[261]);
fa fau_0_262(a_i_c[262],a_i_s[262],b_i_c[262],c_t[262],s_t[262]);
fa fau_0_263(a_i_c[263],a_i_s[263],b_i_c[263],c_t[263],s_t[263]);
fa fau_0_264(a_i_c[264],a_i_s[264],b_i_c[264],c_t[264],s_t[264]);
fa fau_0_265(a_i_c[265],a_i_s[265],b_i_c[265],c_t[265],s_t[265]);
fa fau_0_266(a_i_c[266],a_i_s[266],b_i_c[266],c_t[266],s_t[266]);
fa fau_0_267(a_i_c[267],a_i_s[267],b_i_c[267],c_t[267],s_t[267]);
fa fau_0_268(a_i_c[268],a_i_s[268],b_i_c[268],c_t[268],s_t[268]);
fa fau_0_269(a_i_c[269],a_i_s[269],b_i_c[269],c_t[269],s_t[269]);
fa fau_0_270(a_i_c[270],a_i_s[270],b_i_c[270],c_t[270],s_t[270]);
fa fau_0_271(a_i_c[271],a_i_s[271],b_i_c[271],c_t[271],s_t[271]);
fa fau_0_272(a_i_c[272],a_i_s[272],b_i_c[272],c_t[272],s_t[272]);
fa fau_0_273(a_i_c[273],a_i_s[273],b_i_c[273],c_t[273],s_t[273]);
fa fau_0_274(a_i_c[274],a_i_s[274],b_i_c[274],c_t[274],s_t[274]);
fa fau_0_275(a_i_c[275],a_i_s[275],b_i_c[275],c_t[275],s_t[275]);
fa fau_0_276(a_i_c[276],a_i_s[276],b_i_c[276],c_t[276],s_t[276]);
fa fau_0_277(a_i_c[277],a_i_s[277],b_i_c[277],c_t[277],s_t[277]);
fa fau_0_278(a_i_c[278],a_i_s[278],b_i_c[278],c_t[278],s_t[278]);
fa fau_0_279(a_i_c[279],a_i_s[279],b_i_c[279],c_t[279],s_t[279]);
fa fau_0_280(a_i_c[280],a_i_s[280],b_i_c[280],c_t[280],s_t[280]);
fa fau_0_281(a_i_c[281],a_i_s[281],b_i_c[281],c_t[281],s_t[281]);
fa fau_0_282(a_i_c[282],a_i_s[282],b_i_c[282],c_t[282],s_t[282]);
fa fau_0_283(a_i_c[283],a_i_s[283],b_i_c[283],c_t[283],s_t[283]);
fa fau_0_284(a_i_c[284],a_i_s[284],b_i_c[284],c_t[284],s_t[284]);
fa fau_0_285(a_i_c[285],a_i_s[285],b_i_c[285],c_t[285],s_t[285]);
fa fau_0_286(a_i_c[286],a_i_s[286],b_i_c[286],c_t[286],s_t[286]);
fa fau_0_287(a_i_c[287],a_i_s[287],b_i_c[287],c_t[287],s_t[287]);
fa fau_0_288(a_i_c[288],a_i_s[288],b_i_c[288],c_t[288],s_t[288]);
fa fau_0_289(a_i_c[289],a_i_s[289],b_i_c[289],c_t[289],s_t[289]);
fa fau_0_290(a_i_c[290],a_i_s[290],b_i_c[290],c_t[290],s_t[290]);
fa fau_0_291(a_i_c[291],a_i_s[291],b_i_c[291],c_t[291],s_t[291]);
fa fau_0_292(a_i_c[292],a_i_s[292],b_i_c[292],c_t[292],s_t[292]);
fa fau_0_293(a_i_c[293],a_i_s[293],b_i_c[293],c_t[293],s_t[293]);
fa fau_0_294(a_i_c[294],a_i_s[294],b_i_c[294],c_t[294],s_t[294]);
fa fau_0_295(a_i_c[295],a_i_s[295],b_i_c[295],c_t[295],s_t[295]);
fa fau_0_296(a_i_c[296],a_i_s[296],b_i_c[296],c_t[296],s_t[296]);
fa fau_0_297(a_i_c[297],a_i_s[297],b_i_c[297],c_t[297],s_t[297]);
fa fau_0_298(a_i_c[298],a_i_s[298],b_i_c[298],c_t[298],s_t[298]);
fa fau_0_299(a_i_c[299],a_i_s[299],b_i_c[299],c_t[299],s_t[299]);
fa fau_0_300(a_i_c[300],a_i_s[300],b_i_c[300],c_t[300],s_t[300]);
fa fau_0_301(a_i_c[301],a_i_s[301],b_i_c[301],c_t[301],s_t[301]);
fa fau_0_302(a_i_c[302],a_i_s[302],b_i_c[302],c_t[302],s_t[302]);
fa fau_0_303(a_i_c[303],a_i_s[303],b_i_c[303],c_t[303],s_t[303]);
fa fau_0_304(a_i_c[304],a_i_s[304],b_i_c[304],c_t[304],s_t[304]);
fa fau_0_305(a_i_c[305],a_i_s[305],b_i_c[305],c_t[305],s_t[305]);
fa fau_0_306(a_i_c[306],a_i_s[306],b_i_c[306],c_t[306],s_t[306]);
fa fau_0_307(a_i_c[307],a_i_s[307],b_i_c[307],c_t[307],s_t[307]);
fa fau_0_308(a_i_c[308],a_i_s[308],b_i_c[308],c_t[308],s_t[308]);
fa fau_0_309(a_i_c[309],a_i_s[309],b_i_c[309],c_t[309],s_t[309]);
fa fau_0_310(a_i_c[310],a_i_s[310],b_i_c[310],c_t[310],s_t[310]);
fa fau_0_311(a_i_c[311],a_i_s[311],b_i_c[311],c_t[311],s_t[311]);
fa fau_0_312(a_i_c[312],a_i_s[312],b_i_c[312],c_t[312],s_t[312]);
fa fau_0_313(a_i_c[313],a_i_s[313],b_i_c[313],c_t[313],s_t[313]);
fa fau_0_314(a_i_c[314],a_i_s[314],b_i_c[314],c_t[314],s_t[314]);
fa fau_0_315(a_i_c[315],a_i_s[315],b_i_c[315],c_t[315],s_t[315]);
fa fau_0_316(a_i_c[316],a_i_s[316],b_i_c[316],c_t[316],s_t[316]);
fa fau_0_317(a_i_c[317],a_i_s[317],b_i_c[317],c_t[317],s_t[317]);
fa fau_0_318(a_i_c[318],a_i_s[318],b_i_c[318],c_t[318],s_t[318]);
fa fau_0_319(a_i_c[319],a_i_s[319],b_i_c[319],c_t[319],s_t[319]);
fa fau_0_320(a_i_c[320],a_i_s[320],b_i_c[320],c_t[320],s_t[320]);
fa fau_0_321(a_i_c[321],a_i_s[321],b_i_c[321],c_t[321],s_t[321]);
fa fau_0_322(a_i_c[322],a_i_s[322],b_i_c[322],c_t[322],s_t[322]);
fa fau_0_323(a_i_c[323],a_i_s[323],b_i_c[323],c_t[323],s_t[323]);
fa fau_0_324(a_i_c[324],a_i_s[324],b_i_c[324],c_t[324],s_t[324]);
fa fau_0_325(a_i_c[325],a_i_s[325],b_i_c[325],c_t[325],s_t[325]);
fa fau_0_326(a_i_c[326],a_i_s[326],b_i_c[326],c_t[326],s_t[326]);
fa fau_0_327(a_i_c[327],a_i_s[327],b_i_c[327],c_t[327],s_t[327]);
fa fau_0_328(a_i_c[328],a_i_s[328],b_i_c[328],c_t[328],s_t[328]);
fa fau_0_329(a_i_c[329],a_i_s[329],b_i_c[329],c_t[329],s_t[329]);
fa fau_0_330(a_i_c[330],a_i_s[330],b_i_c[330],c_t[330],s_t[330]);
fa fau_0_331(a_i_c[331],a_i_s[331],b_i_c[331],c_t[331],s_t[331]);
fa fau_0_332(a_i_c[332],a_i_s[332],b_i_c[332],c_t[332],s_t[332]);
fa fau_0_333(a_i_c[333],a_i_s[333],b_i_c[333],c_t[333],s_t[333]);
fa fau_0_334(a_i_c[334],a_i_s[334],b_i_c[334],c_t[334],s_t[334]);
fa fau_0_335(a_i_c[335],a_i_s[335],b_i_c[335],c_t[335],s_t[335]);
fa fau_0_336(a_i_c[336],a_i_s[336],b_i_c[336],c_t[336],s_t[336]);
fa fau_0_337(a_i_c[337],a_i_s[337],b_i_c[337],c_t[337],s_t[337]);
fa fau_0_338(a_i_c[338],a_i_s[338],b_i_c[338],c_t[338],s_t[338]);
fa fau_0_339(a_i_c[339],a_i_s[339],b_i_c[339],c_t[339],s_t[339]);
fa fau_0_340(a_i_c[340],a_i_s[340],b_i_c[340],c_t[340],s_t[340]);
fa fau_0_341(a_i_c[341],a_i_s[341],b_i_c[341],c_t[341],s_t[341]);
fa fau_0_342(a_i_c[342],a_i_s[342],b_i_c[342],c_t[342],s_t[342]);
fa fau_0_343(a_i_c[343],a_i_s[343],b_i_c[343],c_t[343],s_t[343]);
fa fau_0_344(a_i_c[344],a_i_s[344],b_i_c[344],c_t[344],s_t[344]);
fa fau_0_345(a_i_c[345],a_i_s[345],b_i_c[345],c_t[345],s_t[345]);
fa fau_0_346(a_i_c[346],a_i_s[346],b_i_c[346],c_t[346],s_t[346]);
fa fau_0_347(a_i_c[347],a_i_s[347],b_i_c[347],c_t[347],s_t[347]);
fa fau_0_348(a_i_c[348],a_i_s[348],b_i_c[348],c_t[348],s_t[348]);
fa fau_0_349(a_i_c[349],a_i_s[349],b_i_c[349],c_t[349],s_t[349]);
fa fau_0_350(a_i_c[350],a_i_s[350],b_i_c[350],c_t[350],s_t[350]);
fa fau_0_351(a_i_c[351],a_i_s[351],b_i_c[351],c_t[351],s_t[351]);
fa fau_0_352(a_i_c[352],a_i_s[352],b_i_c[352],c_t[352],s_t[352]);
fa fau_0_353(a_i_c[353],a_i_s[353],b_i_c[353],c_t[353],s_t[353]);
fa fau_0_354(a_i_c[354],a_i_s[354],b_i_c[354],c_t[354],s_t[354]);
fa fau_0_355(a_i_c[355],a_i_s[355],b_i_c[355],c_t[355],s_t[355]);
fa fau_0_356(a_i_c[356],a_i_s[356],b_i_c[356],c_t[356],s_t[356]);
fa fau_0_357(a_i_c[357],a_i_s[357],b_i_c[357],c_t[357],s_t[357]);
fa fau_0_358(a_i_c[358],a_i_s[358],b_i_c[358],c_t[358],s_t[358]);
fa fau_0_359(a_i_c[359],a_i_s[359],b_i_c[359],c_t[359],s_t[359]);
fa fau_0_360(a_i_c[360],a_i_s[360],b_i_c[360],c_t[360],s_t[360]);
fa fau_0_361(a_i_c[361],a_i_s[361],b_i_c[361],c_t[361],s_t[361]);
fa fau_0_362(a_i_c[362],a_i_s[362],b_i_c[362],c_t[362],s_t[362]);
fa fau_0_363(a_i_c[363],a_i_s[363],b_i_c[363],c_t[363],s_t[363]);
fa fau_0_364(a_i_c[364],a_i_s[364],b_i_c[364],c_t[364],s_t[364]);
fa fau_0_365(a_i_c[365],a_i_s[365],b_i_c[365],c_t[365],s_t[365]);
fa fau_0_366(a_i_c[366],a_i_s[366],b_i_c[366],c_t[366],s_t[366]);
fa fau_0_367(a_i_c[367],a_i_s[367],b_i_c[367],c_t[367],s_t[367]);
fa fau_0_368(a_i_c[368],a_i_s[368],b_i_c[368],c_t[368],s_t[368]);
fa fau_0_369(a_i_c[369],a_i_s[369],b_i_c[369],c_t[369],s_t[369]);
fa fau_0_370(a_i_c[370],a_i_s[370],b_i_c[370],c_t[370],s_t[370]);
fa fau_0_371(a_i_c[371],a_i_s[371],b_i_c[371],c_t[371],s_t[371]);
fa fau_0_372(a_i_c[372],a_i_s[372],b_i_c[372],c_t[372],s_t[372]);
fa fau_0_373(a_i_c[373],a_i_s[373],b_i_c[373],c_t[373],s_t[373]);
fa fau_0_374(a_i_c[374],a_i_s[374],b_i_c[374],c_t[374],s_t[374]);
fa fau_0_375(a_i_c[375],a_i_s[375],b_i_c[375],c_t[375],s_t[375]);
fa fau_0_376(a_i_c[376],a_i_s[376],b_i_c[376],c_t[376],s_t[376]);
fa fau_0_377(a_i_c[377],a_i_s[377],b_i_c[377],c_t[377],s_t[377]);
fa fau_0_378(a_i_c[378],a_i_s[378],b_i_c[378],c_t[378],s_t[378]);
fa fau_0_379(a_i_c[379],a_i_s[379],b_i_c[379],c_t[379],s_t[379]);
fa fau_0_380(a_i_c[380],a_i_s[380],b_i_c[380],c_t[380],s_t[380]);
fa fau_0_381(a_i_c[381],a_i_s[381],b_i_c[381],c_t[381],s_t[381]);
fa fau_0_382(a_i_c[382],a_i_s[382],b_i_c[382],c_t[382],s_t[382]);
fa fau_0_383(a_i_c[383],a_i_s[383],b_i_c[383],c_t[383],s_t[383]);
fa fau_0_384(a_i_c[384],a_i_s[384],b_i_c[384],c_t[384],s_t[384]);
fa fau_0_385(a_i_c[385],a_i_s[385],b_i_c[385],c_t[385],s_t[385]);
fa fau_0_386(a_i_c[386],a_i_s[386],b_i_c[386],c_t[386],s_t[386]);
fa fau_0_387(a_i_c[387],a_i_s[387],b_i_c[387],c_t[387],s_t[387]);
fa fau_0_388(a_i_c[388],a_i_s[388],b_i_c[388],c_t[388],s_t[388]);
fa fau_0_389(a_i_c[389],a_i_s[389],b_i_c[389],c_t[389],s_t[389]);
fa fau_0_390(a_i_c[390],a_i_s[390],b_i_c[390],c_t[390],s_t[390]);
fa fau_0_391(a_i_c[391],a_i_s[391],b_i_c[391],c_t[391],s_t[391]);
fa fau_0_392(a_i_c[392],a_i_s[392],b_i_c[392],c_t[392],s_t[392]);
fa fau_0_393(a_i_c[393],a_i_s[393],b_i_c[393],c_t[393],s_t[393]);
fa fau_0_394(a_i_c[394],a_i_s[394],b_i_c[394],c_t[394],s_t[394]);
fa fau_0_395(a_i_c[395],a_i_s[395],b_i_c[395],c_t[395],s_t[395]);
fa fau_0_396(a_i_c[396],a_i_s[396],b_i_c[396],c_t[396],s_t[396]);
fa fau_0_397(a_i_c[397],a_i_s[397],b_i_c[397],c_t[397],s_t[397]);
fa fau_0_398(a_i_c[398],a_i_s[398],b_i_c[398],c_t[398],s_t[398]);
fa fau_0_399(a_i_c[399],a_i_s[399],b_i_c[399],c_t[399],s_t[399]);
fa fau_0_400(a_i_c[400],a_i_s[400],b_i_c[400],c_t[400],s_t[400]);
fa fau_0_401(a_i_c[401],a_i_s[401],b_i_c[401],c_t[401],s_t[401]);
fa fau_0_402(a_i_c[402],a_i_s[402],b_i_c[402],c_t[402],s_t[402]);
fa fau_0_403(a_i_c[403],a_i_s[403],b_i_c[403],c_t[403],s_t[403]);
fa fau_0_404(a_i_c[404],a_i_s[404],b_i_c[404],c_t[404],s_t[404]);
fa fau_0_405(a_i_c[405],a_i_s[405],b_i_c[405],c_t[405],s_t[405]);
fa fau_0_406(a_i_c[406],a_i_s[406],b_i_c[406],c_t[406],s_t[406]);
fa fau_0_407(a_i_c[407],a_i_s[407],b_i_c[407],c_t[407],s_t[407]);
fa fau_0_408(a_i_c[408],a_i_s[408],b_i_c[408],c_t[408],s_t[408]);
fa fau_0_409(a_i_c[409],a_i_s[409],b_i_c[409],c_t[409],s_t[409]);
fa fau_0_410(a_i_c[410],a_i_s[410],b_i_c[410],c_t[410],s_t[410]);
fa fau_0_411(a_i_c[411],a_i_s[411],b_i_c[411],c_t[411],s_t[411]);
fa fau_0_412(a_i_c[412],a_i_s[412],b_i_c[412],c_t[412],s_t[412]);
fa fau_0_413(a_i_c[413],a_i_s[413],b_i_c[413],c_t[413],s_t[413]);
fa fau_0_414(a_i_c[414],a_i_s[414],b_i_c[414],c_t[414],s_t[414]);
fa fau_0_415(a_i_c[415],a_i_s[415],b_i_c[415],c_t[415],s_t[415]);
fa fau_0_416(a_i_c[416],a_i_s[416],b_i_c[416],c_t[416],s_t[416]);
fa fau_0_417(a_i_c[417],a_i_s[417],b_i_c[417],c_t[417],s_t[417]);
fa fau_0_418(a_i_c[418],a_i_s[418],b_i_c[418],c_t[418],s_t[418]);
fa fau_0_419(a_i_c[419],a_i_s[419],b_i_c[419],c_t[419],s_t[419]);
fa fau_0_420(a_i_c[420],a_i_s[420],b_i_c[420],c_t[420],s_t[420]);
fa fau_0_421(a_i_c[421],a_i_s[421],b_i_c[421],c_t[421],s_t[421]);
fa fau_0_422(a_i_c[422],a_i_s[422],b_i_c[422],c_t[422],s_t[422]);
fa fau_0_423(a_i_c[423],a_i_s[423],b_i_c[423],c_t[423],s_t[423]);
fa fau_0_424(a_i_c[424],a_i_s[424],b_i_c[424],c_t[424],s_t[424]);
fa fau_0_425(a_i_c[425],a_i_s[425],b_i_c[425],c_t[425],s_t[425]);
fa fau_0_426(a_i_c[426],a_i_s[426],b_i_c[426],c_t[426],s_t[426]);
fa fau_0_427(a_i_c[427],a_i_s[427],b_i_c[427],c_t[427],s_t[427]);
fa fau_0_428(a_i_c[428],a_i_s[428],b_i_c[428],c_t[428],s_t[428]);
fa fau_0_429(a_i_c[429],a_i_s[429],b_i_c[429],c_t[429],s_t[429]);
fa fau_0_430(a_i_c[430],a_i_s[430],b_i_c[430],c_t[430],s_t[430]);
fa fau_0_431(a_i_c[431],a_i_s[431],b_i_c[431],c_t[431],s_t[431]);
fa fau_0_432(a_i_c[432],a_i_s[432],b_i_c[432],c_t[432],s_t[432]);
fa fau_0_433(a_i_c[433],a_i_s[433],b_i_c[433],c_t[433],s_t[433]);
fa fau_0_434(a_i_c[434],a_i_s[434],b_i_c[434],c_t[434],s_t[434]);
fa fau_0_435(a_i_c[435],a_i_s[435],b_i_c[435],c_t[435],s_t[435]);
fa fau_0_436(a_i_c[436],a_i_s[436],b_i_c[436],c_t[436],s_t[436]);
fa fau_0_437(a_i_c[437],a_i_s[437],b_i_c[437],c_t[437],s_t[437]);
fa fau_0_438(a_i_c[438],a_i_s[438],b_i_c[438],c_t[438],s_t[438]);
fa fau_0_439(a_i_c[439],a_i_s[439],b_i_c[439],c_t[439],s_t[439]);
fa fau_0_440(a_i_c[440],a_i_s[440],b_i_c[440],c_t[440],s_t[440]);
fa fau_0_441(a_i_c[441],a_i_s[441],b_i_c[441],c_t[441],s_t[441]);
fa fau_0_442(a_i_c[442],a_i_s[442],b_i_c[442],c_t[442],s_t[442]);
fa fau_0_443(a_i_c[443],a_i_s[443],b_i_c[443],c_t[443],s_t[443]);
fa fau_0_444(a_i_c[444],a_i_s[444],b_i_c[444],c_t[444],s_t[444]);
fa fau_0_445(a_i_c[445],a_i_s[445],b_i_c[445],c_t[445],s_t[445]);
fa fau_0_446(a_i_c[446],a_i_s[446],b_i_c[446],c_t[446],s_t[446]);
fa fau_0_447(a_i_c[447],a_i_s[447],b_i_c[447],c_t[447],s_t[447]);
fa fau_0_448(a_i_c[448],a_i_s[448],b_i_c[448],c_t[448],s_t[448]);
fa fau_0_449(a_i_c[449],a_i_s[449],b_i_c[449],c_t[449],s_t[449]);
fa fau_0_450(a_i_c[450],a_i_s[450],b_i_c[450],c_t[450],s_t[450]);
fa fau_0_451(a_i_c[451],a_i_s[451],b_i_c[451],c_t[451],s_t[451]);
fa fau_0_452(a_i_c[452],a_i_s[452],b_i_c[452],c_t[452],s_t[452]);
fa fau_0_453(a_i_c[453],a_i_s[453],b_i_c[453],c_t[453],s_t[453]);
fa fau_0_454(a_i_c[454],a_i_s[454],b_i_c[454],c_t[454],s_t[454]);
fa fau_0_455(a_i_c[455],a_i_s[455],b_i_c[455],c_t[455],s_t[455]);
fa fau_0_456(a_i_c[456],a_i_s[456],b_i_c[456],c_t[456],s_t[456]);
fa fau_0_457(a_i_c[457],a_i_s[457],b_i_c[457],c_t[457],s_t[457]);
fa fau_0_458(a_i_c[458],a_i_s[458],b_i_c[458],c_t[458],s_t[458]);
fa fau_0_459(a_i_c[459],a_i_s[459],b_i_c[459],c_t[459],s_t[459]);
fa fau_0_460(a_i_c[460],a_i_s[460],b_i_c[460],c_t[460],s_t[460]);
fa fau_0_461(a_i_c[461],a_i_s[461],b_i_c[461],c_t[461],s_t[461]);
fa fau_0_462(a_i_c[462],a_i_s[462],b_i_c[462],c_t[462],s_t[462]);
fa fau_0_463(a_i_c[463],a_i_s[463],b_i_c[463],c_t[463],s_t[463]);
fa fau_0_464(a_i_c[464],a_i_s[464],b_i_c[464],c_t[464],s_t[464]);
fa fau_0_465(a_i_c[465],a_i_s[465],b_i_c[465],c_t[465],s_t[465]);
fa fau_0_466(a_i_c[466],a_i_s[466],b_i_c[466],c_t[466],s_t[466]);
fa fau_0_467(a_i_c[467],a_i_s[467],b_i_c[467],c_t[467],s_t[467]);
fa fau_0_468(a_i_c[468],a_i_s[468],b_i_c[468],c_t[468],s_t[468]);
fa fau_0_469(a_i_c[469],a_i_s[469],b_i_c[469],c_t[469],s_t[469]);
fa fau_0_470(a_i_c[470],a_i_s[470],b_i_c[470],c_t[470],s_t[470]);
fa fau_0_471(a_i_c[471],a_i_s[471],b_i_c[471],c_t[471],s_t[471]);
fa fau_0_472(a_i_c[472],a_i_s[472],b_i_c[472],c_t[472],s_t[472]);
fa fau_0_473(a_i_c[473],a_i_s[473],b_i_c[473],c_t[473],s_t[473]);
fa fau_0_474(a_i_c[474],a_i_s[474],b_i_c[474],c_t[474],s_t[474]);
fa fau_0_475(a_i_c[475],a_i_s[475],b_i_c[475],c_t[475],s_t[475]);
fa fau_0_476(a_i_c[476],a_i_s[476],b_i_c[476],c_t[476],s_t[476]);
fa fau_0_477(a_i_c[477],a_i_s[477],b_i_c[477],c_t[477],s_t[477]);
fa fau_0_478(a_i_c[478],a_i_s[478],b_i_c[478],c_t[478],s_t[478]);
fa fau_0_479(a_i_c[479],a_i_s[479],b_i_c[479],c_t[479],s_t[479]);
fa fau_0_480(a_i_c[480],a_i_s[480],b_i_c[480],c_t[480],s_t[480]);
fa fau_0_481(a_i_c[481],a_i_s[481],b_i_c[481],c_t[481],s_t[481]);
fa fau_0_482(a_i_c[482],a_i_s[482],b_i_c[482],c_t[482],s_t[482]);
fa fau_0_483(a_i_c[483],a_i_s[483],b_i_c[483],c_t[483],s_t[483]);
fa fau_0_484(a_i_c[484],a_i_s[484],b_i_c[484],c_t[484],s_t[484]);
fa fau_0_485(a_i_c[485],a_i_s[485],b_i_c[485],c_t[485],s_t[485]);
fa fau_0_486(a_i_c[486],a_i_s[486],b_i_c[486],c_t[486],s_t[486]);
fa fau_0_487(a_i_c[487],a_i_s[487],b_i_c[487],c_t[487],s_t[487]);
fa fau_0_488(a_i_c[488],a_i_s[488],b_i_c[488],c_t[488],s_t[488]);
fa fau_0_489(a_i_c[489],a_i_s[489],b_i_c[489],c_t[489],s_t[489]);
fa fau_0_490(a_i_c[490],a_i_s[490],b_i_c[490],c_t[490],s_t[490]);
fa fau_0_491(a_i_c[491],a_i_s[491],b_i_c[491],c_t[491],s_t[491]);
fa fau_0_492(a_i_c[492],a_i_s[492],b_i_c[492],c_t[492],s_t[492]);
fa fau_0_493(a_i_c[493],a_i_s[493],b_i_c[493],c_t[493],s_t[493]);
fa fau_0_494(a_i_c[494],a_i_s[494],b_i_c[494],c_t[494],s_t[494]);
fa fau_0_495(a_i_c[495],a_i_s[495],b_i_c[495],c_t[495],s_t[495]);
fa fau_0_496(a_i_c[496],a_i_s[496],b_i_c[496],c_t[496],s_t[496]);
fa fau_0_497(a_i_c[497],a_i_s[497],b_i_c[497],c_t[497],s_t[497]);
fa fau_0_498(a_i_c[498],a_i_s[498],b_i_c[498],c_t[498],s_t[498]);
fa fau_0_499(a_i_c[499],a_i_s[499],b_i_c[499],c_t[499],s_t[499]);
fa fau_0_500(a_i_c[500],a_i_s[500],b_i_c[500],c_t[500],s_t[500]);
fa fau_0_501(a_i_c[501],a_i_s[501],b_i_c[501],c_t[501],s_t[501]);
fa fau_0_502(a_i_c[502],a_i_s[502],b_i_c[502],c_t[502],s_t[502]);
fa fau_0_503(a_i_c[503],a_i_s[503],b_i_c[503],c_t[503],s_t[503]);
fa fau_0_504(a_i_c[504],a_i_s[504],b_i_c[504],c_t[504],s_t[504]);
fa fau_0_505(a_i_c[505],a_i_s[505],b_i_c[505],c_t[505],s_t[505]);
fa fau_0_506(a_i_c[506],a_i_s[506],b_i_c[506],c_t[506],s_t[506]);
fa fau_0_507(a_i_c[507],a_i_s[507],b_i_c[507],c_t[507],s_t[507]);
fa fau_0_508(a_i_c[508],a_i_s[508],b_i_c[508],c_t[508],s_t[508]);
fa fau_0_509(a_i_c[509],a_i_s[509],b_i_c[509],c_t[509],s_t[509]);
fa fau_0_510(a_i_c[510],a_i_s[510],b_i_c[510],c_t[510],s_t[510]);
fa fau_0_511(a_i_c[511],a_i_s[511],b_i_c[511],c_t[511],s_t[511]);
fa fau_0_512(a_i_c[512],a_i_s[512],b_i_c[512],c_t[512],s_t[512]);
fa fau_0_513(a_i_c[513],a_i_s[513],b_i_c[513],c_t[513],s_t[513]);
fa fau_0_514(a_i_c[514],a_i_s[514],b_i_c[514],c_t[514],s_t[514]);
fa fau_0_515(a_i_c[515],a_i_s[515],b_i_c[515],c_t[515],s_t[515]);
fa fau_0_516(a_i_c[516],a_i_s[516],b_i_c[516],c_t[516],s_t[516]);
fa fau_0_517(a_i_c[517],a_i_s[517],b_i_c[517],c_t[517],s_t[517]);
fa fau_0_518(a_i_c[518],a_i_s[518],b_i_c[518],c_t[518],s_t[518]);
fa fau_0_519(a_i_c[519],a_i_s[519],b_i_c[519],c_t[519],s_t[519]);
fa fau_0_520(a_i_c[520],a_i_s[520],b_i_c[520],c_t[520],s_t[520]);
fa fau_0_521(a_i_c[521],a_i_s[521],b_i_c[521],c_t[521],s_t[521]);
fa fau_0_522(a_i_c[522],a_i_s[522],b_i_c[522],c_t[522],s_t[522]);
fa fau_0_523(a_i_c[523],a_i_s[523],b_i_c[523],c_t[523],s_t[523]);
fa fau_0_524(a_i_c[524],a_i_s[524],b_i_c[524],c_t[524],s_t[524]);
fa fau_0_525(a_i_c[525],a_i_s[525],b_i_c[525],c_t[525],s_t[525]);
fa fau_0_526(a_i_c[526],a_i_s[526],b_i_c[526],c_t[526],s_t[526]);
fa fau_0_527(a_i_c[527],a_i_s[527],b_i_c[527],c_t[527],s_t[527]);
fa fau_0_528(a_i_c[528],a_i_s[528],b_i_c[528],c_t[528],s_t[528]);
fa fau_0_529(a_i_c[529],a_i_s[529],b_i_c[529],c_t[529],s_t[529]);
fa fau_0_530(a_i_c[530],a_i_s[530],b_i_c[530],c_t[530],s_t[530]);
fa fau_0_531(a_i_c[531],a_i_s[531],b_i_c[531],c_t[531],s_t[531]);
fa fau_0_532(a_i_c[532],a_i_s[532],b_i_c[532],c_t[532],s_t[532]);
fa fau_0_533(a_i_c[533],a_i_s[533],b_i_c[533],c_t[533],s_t[533]);
fa fau_0_534(a_i_c[534],a_i_s[534],b_i_c[534],c_t[534],s_t[534]);
fa fau_0_535(a_i_c[535],a_i_s[535],b_i_c[535],c_t[535],s_t[535]);
fa fau_0_536(a_i_c[536],a_i_s[536],b_i_c[536],c_t[536],s_t[536]);
fa fau_0_537(a_i_c[537],a_i_s[537],b_i_c[537],c_t[537],s_t[537]);
fa fau_0_538(a_i_c[538],a_i_s[538],b_i_c[538],c_t[538],s_t[538]);
fa fau_0_539(a_i_c[539],a_i_s[539],b_i_c[539],c_t[539],s_t[539]);
fa fau_0_540(a_i_c[540],a_i_s[540],b_i_c[540],c_t[540],s_t[540]);
fa fau_0_541(a_i_c[541],a_i_s[541],b_i_c[541],c_t[541],s_t[541]);
fa fau_0_542(a_i_c[542],a_i_s[542],b_i_c[542],c_t[542],s_t[542]);
fa fau_0_543(a_i_c[543],a_i_s[543],b_i_c[543],c_t[543],s_t[543]);
fa fau_0_544(a_i_c[544],a_i_s[544],b_i_c[544],c_t[544],s_t[544]);
fa fau_0_545(a_i_c[545],a_i_s[545],b_i_c[545],c_t[545],s_t[545]);
fa fau_0_546(a_i_c[546],a_i_s[546],b_i_c[546],c_t[546],s_t[546]);
fa fau_0_547(a_i_c[547],a_i_s[547],b_i_c[547],c_t[547],s_t[547]);
fa fau_0_548(a_i_c[548],a_i_s[548],b_i_c[548],c_t[548],s_t[548]);
fa fau_0_549(a_i_c[549],a_i_s[549],b_i_c[549],c_t[549],s_t[549]);
fa fau_0_550(a_i_c[550],a_i_s[550],b_i_c[550],c_t[550],s_t[550]);
fa fau_0_551(a_i_c[551],a_i_s[551],b_i_c[551],c_t[551],s_t[551]);
fa fau_0_552(a_i_c[552],a_i_s[552],b_i_c[552],c_t[552],s_t[552]);
fa fau_0_553(a_i_c[553],a_i_s[553],b_i_c[553],c_t[553],s_t[553]);
fa fau_0_554(a_i_c[554],a_i_s[554],b_i_c[554],c_t[554],s_t[554]);
fa fau_0_555(a_i_c[555],a_i_s[555],b_i_c[555],c_t[555],s_t[555]);
fa fau_0_556(a_i_c[556],a_i_s[556],b_i_c[556],c_t[556],s_t[556]);
fa fau_0_557(a_i_c[557],a_i_s[557],b_i_c[557],c_t[557],s_t[557]);
fa fau_0_558(a_i_c[558],a_i_s[558],b_i_c[558],c_t[558],s_t[558]);
fa fau_0_559(a_i_c[559],a_i_s[559],b_i_c[559],c_t[559],s_t[559]);
fa fau_0_560(a_i_c[560],a_i_s[560],b_i_c[560],c_t[560],s_t[560]);
fa fau_0_561(a_i_c[561],a_i_s[561],b_i_c[561],c_t[561],s_t[561]);
fa fau_0_562(a_i_c[562],a_i_s[562],b_i_c[562],c_t[562],s_t[562]);
fa fau_0_563(a_i_c[563],a_i_s[563],b_i_c[563],c_t[563],s_t[563]);
fa fau_0_564(a_i_c[564],a_i_s[564],b_i_c[564],c_t[564],s_t[564]);
fa fau_0_565(a_i_c[565],a_i_s[565],b_i_c[565],c_t[565],s_t[565]);
fa fau_0_566(a_i_c[566],a_i_s[566],b_i_c[566],c_t[566],s_t[566]);
fa fau_0_567(a_i_c[567],a_i_s[567],b_i_c[567],c_t[567],s_t[567]);
fa fau_0_568(a_i_c[568],a_i_s[568],b_i_c[568],c_t[568],s_t[568]);
fa fau_0_569(a_i_c[569],a_i_s[569],b_i_c[569],c_t[569],s_t[569]);
fa fau_0_570(a_i_c[570],a_i_s[570],b_i_c[570],c_t[570],s_t[570]);
fa fau_0_571(a_i_c[571],a_i_s[571],b_i_c[571],c_t[571],s_t[571]);
fa fau_0_572(a_i_c[572],a_i_s[572],b_i_c[572],c_t[572],s_t[572]);
fa fau_0_573(a_i_c[573],a_i_s[573],b_i_c[573],c_t[573],s_t[573]);
fa fau_0_574(a_i_c[574],a_i_s[574],b_i_c[574],c_t[574],s_t[574]);
fa fau_0_575(a_i_c[575],a_i_s[575],b_i_c[575],c_t[575],s_t[575]);
fa fau_0_576(a_i_c[576],a_i_s[576],b_i_c[576],c_t[576],s_t[576]);
fa fau_0_577(a_i_c[577],a_i_s[577],b_i_c[577],c_t[577],s_t[577]);
fa fau_0_578(a_i_c[578],a_i_s[578],b_i_c[578],c_t[578],s_t[578]);
fa fau_0_579(a_i_c[579],a_i_s[579],b_i_c[579],c_t[579],s_t[579]);
fa fau_0_580(a_i_c[580],a_i_s[580],b_i_c[580],c_t[580],s_t[580]);
fa fau_0_581(a_i_c[581],a_i_s[581],b_i_c[581],c_t[581],s_t[581]);
fa fau_0_582(a_i_c[582],a_i_s[582],b_i_c[582],c_t[582],s_t[582]);
fa fau_0_583(a_i_c[583],a_i_s[583],b_i_c[583],c_t[583],s_t[583]);
fa fau_0_584(a_i_c[584],a_i_s[584],b_i_c[584],c_t[584],s_t[584]);
fa fau_0_585(a_i_c[585],a_i_s[585],b_i_c[585],c_t[585],s_t[585]);
fa fau_0_586(a_i_c[586],a_i_s[586],b_i_c[586],c_t[586],s_t[586]);
fa fau_0_587(a_i_c[587],a_i_s[587],b_i_c[587],c_t[587],s_t[587]);
fa fau_0_588(a_i_c[588],a_i_s[588],b_i_c[588],c_t[588],s_t[588]);
fa fau_0_589(a_i_c[589],a_i_s[589],b_i_c[589],c_t[589],s_t[589]);
fa fau_0_590(a_i_c[590],a_i_s[590],b_i_c[590],c_t[590],s_t[590]);
fa fau_0_591(a_i_c[591],a_i_s[591],b_i_c[591],c_t[591],s_t[591]);
fa fau_0_592(a_i_c[592],a_i_s[592],b_i_c[592],c_t[592],s_t[592]);
fa fau_0_593(a_i_c[593],a_i_s[593],b_i_c[593],c_t[593],s_t[593]);
fa fau_0_594(a_i_c[594],a_i_s[594],b_i_c[594],c_t[594],s_t[594]);
fa fau_0_595(a_i_c[595],a_i_s[595],b_i_c[595],c_t[595],s_t[595]);
fa fau_0_596(a_i_c[596],a_i_s[596],b_i_c[596],c_t[596],s_t[596]);
fa fau_0_597(a_i_c[597],a_i_s[597],b_i_c[597],c_t[597],s_t[597]);
fa fau_0_598(a_i_c[598],a_i_s[598],b_i_c[598],c_t[598],s_t[598]);
fa fau_0_599(a_i_c[599],a_i_s[599],b_i_c[599],c_t[599],s_t[599]);
fa fau_0_600(a_i_c[600],a_i_s[600],b_i_c[600],c_t[600],s_t[600]);
fa fau_0_601(a_i_c[601],a_i_s[601],b_i_c[601],c_t[601],s_t[601]);
fa fau_0_602(a_i_c[602],a_i_s[602],b_i_c[602],c_t[602],s_t[602]);
fa fau_0_603(a_i_c[603],a_i_s[603],b_i_c[603],c_t[603],s_t[603]);
fa fau_0_604(a_i_c[604],a_i_s[604],b_i_c[604],c_t[604],s_t[604]);
fa fau_0_605(a_i_c[605],a_i_s[605],b_i_c[605],c_t[605],s_t[605]);
fa fau_0_606(a_i_c[606],a_i_s[606],b_i_c[606],c_t[606],s_t[606]);
fa fau_0_607(a_i_c[607],a_i_s[607],b_i_c[607],c_t[607],s_t[607]);
fa fau_0_608(a_i_c[608],a_i_s[608],b_i_c[608],c_t[608],s_t[608]);
fa fau_0_609(a_i_c[609],a_i_s[609],b_i_c[609],c_t[609],s_t[609]);
fa fau_0_610(a_i_c[610],a_i_s[610],b_i_c[610],c_t[610],s_t[610]);
fa fau_0_611(a_i_c[611],a_i_s[611],b_i_c[611],c_t[611],s_t[611]);
fa fau_0_612(a_i_c[612],a_i_s[612],b_i_c[612],c_t[612],s_t[612]);
fa fau_0_613(a_i_c[613],a_i_s[613],b_i_c[613],c_t[613],s_t[613]);
fa fau_0_614(a_i_c[614],a_i_s[614],b_i_c[614],c_t[614],s_t[614]);
fa fau_0_615(a_i_c[615],a_i_s[615],b_i_c[615],c_t[615],s_t[615]);
fa fau_0_616(a_i_c[616],a_i_s[616],b_i_c[616],c_t[616],s_t[616]);
fa fau_0_617(a_i_c[617],a_i_s[617],b_i_c[617],c_t[617],s_t[617]);
fa fau_0_618(a_i_c[618],a_i_s[618],b_i_c[618],c_t[618],s_t[618]);
fa fau_0_619(a_i_c[619],a_i_s[619],b_i_c[619],c_t[619],s_t[619]);
fa fau_0_620(a_i_c[620],a_i_s[620],b_i_c[620],c_t[620],s_t[620]);
fa fau_0_621(a_i_c[621],a_i_s[621],b_i_c[621],c_t[621],s_t[621]);
fa fau_0_622(a_i_c[622],a_i_s[622],b_i_c[622],c_t[622],s_t[622]);
fa fau_0_623(a_i_c[623],a_i_s[623],b_i_c[623],c_t[623],s_t[623]);
fa fau_0_624(a_i_c[624],a_i_s[624],b_i_c[624],c_t[624],s_t[624]);
fa fau_0_625(a_i_c[625],a_i_s[625],b_i_c[625],c_t[625],s_t[625]);
fa fau_0_626(a_i_c[626],a_i_s[626],b_i_c[626],c_t[626],s_t[626]);
fa fau_0_627(a_i_c[627],a_i_s[627],b_i_c[627],c_t[627],s_t[627]);
fa fau_0_628(a_i_c[628],a_i_s[628],b_i_c[628],c_t[628],s_t[628]);
fa fau_0_629(a_i_c[629],a_i_s[629],b_i_c[629],c_t[629],s_t[629]);
fa fau_0_630(a_i_c[630],a_i_s[630],b_i_c[630],c_t[630],s_t[630]);
fa fau_0_631(a_i_c[631],a_i_s[631],b_i_c[631],c_t[631],s_t[631]);
fa fau_0_632(a_i_c[632],a_i_s[632],b_i_c[632],c_t[632],s_t[632]);
fa fau_0_633(a_i_c[633],a_i_s[633],b_i_c[633],c_t[633],s_t[633]);
fa fau_0_634(a_i_c[634],a_i_s[634],b_i_c[634],c_t[634],s_t[634]);
fa fau_0_635(a_i_c[635],a_i_s[635],b_i_c[635],c_t[635],s_t[635]);
fa fau_0_636(a_i_c[636],a_i_s[636],b_i_c[636],c_t[636],s_t[636]);
fa fau_0_637(a_i_c[637],a_i_s[637],b_i_c[637],c_t[637],s_t[637]);
fa fau_0_638(a_i_c[638],a_i_s[638],b_i_c[638],c_t[638],s_t[638]);
fa fau_0_639(a_i_c[639],a_i_s[639],b_i_c[639],c_t[639],s_t[639]);
fa fau_0_640(a_i_c[640],a_i_s[640],b_i_c[640],c_t[640],s_t[640]);
fa fau_0_641(a_i_c[641],a_i_s[641],b_i_c[641],c_t[641],s_t[641]);
fa fau_0_642(a_i_c[642],a_i_s[642],b_i_c[642],c_t[642],s_t[642]);
fa fau_0_643(a_i_c[643],a_i_s[643],b_i_c[643],c_t[643],s_t[643]);
fa fau_0_644(a_i_c[644],a_i_s[644],b_i_c[644],c_t[644],s_t[644]);
fa fau_0_645(a_i_c[645],a_i_s[645],b_i_c[645],c_t[645],s_t[645]);
fa fau_0_646(a_i_c[646],a_i_s[646],b_i_c[646],c_t[646],s_t[646]);
fa fau_0_647(a_i_c[647],a_i_s[647],b_i_c[647],c_t[647],s_t[647]);
fa fau_0_648(a_i_c[648],a_i_s[648],b_i_c[648],c_t[648],s_t[648]);
fa fau_0_649(a_i_c[649],a_i_s[649],b_i_c[649],c_t[649],s_t[649]);
fa fau_0_650(a_i_c[650],a_i_s[650],b_i_c[650],c_t[650],s_t[650]);
fa fau_0_651(a_i_c[651],a_i_s[651],b_i_c[651],c_t[651],s_t[651]);
fa fau_0_652(a_i_c[652],a_i_s[652],b_i_c[652],c_t[652],s_t[652]);
fa fau_0_653(a_i_c[653],a_i_s[653],b_i_c[653],c_t[653],s_t[653]);
fa fau_0_654(a_i_c[654],a_i_s[654],b_i_c[654],c_t[654],s_t[654]);
fa fau_0_655(a_i_c[655],a_i_s[655],b_i_c[655],c_t[655],s_t[655]);
fa fau_0_656(a_i_c[656],a_i_s[656],b_i_c[656],c_t[656],s_t[656]);
fa fau_0_657(a_i_c[657],a_i_s[657],b_i_c[657],c_t[657],s_t[657]);
fa fau_0_658(a_i_c[658],a_i_s[658],b_i_c[658],c_t[658],s_t[658]);
fa fau_0_659(a_i_c[659],a_i_s[659],b_i_c[659],c_t[659],s_t[659]);
fa fau_0_660(a_i_c[660],a_i_s[660],b_i_c[660],c_t[660],s_t[660]);
fa fau_0_661(a_i_c[661],a_i_s[661],b_i_c[661],c_t[661],s_t[661]);
fa fau_0_662(a_i_c[662],a_i_s[662],b_i_c[662],c_t[662],s_t[662]);
fa fau_0_663(a_i_c[663],a_i_s[663],b_i_c[663],c_t[663],s_t[663]);
fa fau_0_664(a_i_c[664],a_i_s[664],b_i_c[664],c_t[664],s_t[664]);
fa fau_0_665(a_i_c[665],a_i_s[665],b_i_c[665],c_t[665],s_t[665]);
fa fau_0_666(a_i_c[666],a_i_s[666],b_i_c[666],c_t[666],s_t[666]);
fa fau_0_667(a_i_c[667],a_i_s[667],b_i_c[667],c_t[667],s_t[667]);
fa fau_0_668(a_i_c[668],a_i_s[668],b_i_c[668],c_t[668],s_t[668]);
fa fau_0_669(a_i_c[669],a_i_s[669],b_i_c[669],c_t[669],s_t[669]);
fa fau_0_670(a_i_c[670],a_i_s[670],b_i_c[670],c_t[670],s_t[670]);
fa fau_0_671(a_i_c[671],a_i_s[671],b_i_c[671],c_t[671],s_t[671]);
fa fau_0_672(a_i_c[672],a_i_s[672],b_i_c[672],c_t[672],s_t[672]);
fa fau_0_673(a_i_c[673],a_i_s[673],b_i_c[673],c_t[673],s_t[673]);
fa fau_0_674(a_i_c[674],a_i_s[674],b_i_c[674],c_t[674],s_t[674]);
fa fau_0_675(a_i_c[675],a_i_s[675],b_i_c[675],c_t[675],s_t[675]);
fa fau_0_676(a_i_c[676],a_i_s[676],b_i_c[676],c_t[676],s_t[676]);
fa fau_0_677(a_i_c[677],a_i_s[677],b_i_c[677],c_t[677],s_t[677]);
fa fau_0_678(a_i_c[678],a_i_s[678],b_i_c[678],c_t[678],s_t[678]);
fa fau_0_679(a_i_c[679],a_i_s[679],b_i_c[679],c_t[679],s_t[679]);
fa fau_0_680(a_i_c[680],a_i_s[680],b_i_c[680],c_t[680],s_t[680]);
fa fau_0_681(a_i_c[681],a_i_s[681],b_i_c[681],c_t[681],s_t[681]);
fa fau_0_682(a_i_c[682],a_i_s[682],b_i_c[682],c_t[682],s_t[682]);
fa fau_0_683(a_i_c[683],a_i_s[683],b_i_c[683],c_t[683],s_t[683]);
fa fau_0_684(a_i_c[684],a_i_s[684],b_i_c[684],c_t[684],s_t[684]);
fa fau_0_685(a_i_c[685],a_i_s[685],b_i_c[685],c_t[685],s_t[685]);
fa fau_0_686(a_i_c[686],a_i_s[686],b_i_c[686],c_t[686],s_t[686]);
fa fau_0_687(a_i_c[687],a_i_s[687],b_i_c[687],c_t[687],s_t[687]);
fa fau_0_688(a_i_c[688],a_i_s[688],b_i_c[688],c_t[688],s_t[688]);
fa fau_0_689(a_i_c[689],a_i_s[689],b_i_c[689],c_t[689],s_t[689]);
fa fau_0_690(a_i_c[690],a_i_s[690],b_i_c[690],c_t[690],s_t[690]);
fa fau_0_691(a_i_c[691],a_i_s[691],b_i_c[691],c_t[691],s_t[691]);
fa fau_0_692(a_i_c[692],a_i_s[692],b_i_c[692],c_t[692],s_t[692]);
fa fau_0_693(a_i_c[693],a_i_s[693],b_i_c[693],c_t[693],s_t[693]);
fa fau_0_694(a_i_c[694],a_i_s[694],b_i_c[694],c_t[694],s_t[694]);
fa fau_0_695(a_i_c[695],a_i_s[695],b_i_c[695],c_t[695],s_t[695]);
fa fau_0_696(a_i_c[696],a_i_s[696],b_i_c[696],c_t[696],s_t[696]);
fa fau_0_697(a_i_c[697],a_i_s[697],b_i_c[697],c_t[697],s_t[697]);
fa fau_0_698(a_i_c[698],a_i_s[698],b_i_c[698],c_t[698],s_t[698]);
fa fau_0_699(a_i_c[699],a_i_s[699],b_i_c[699],c_t[699],s_t[699]);
fa fau_0_700(a_i_c[700],a_i_s[700],b_i_c[700],c_t[700],s_t[700]);
fa fau_0_701(a_i_c[701],a_i_s[701],b_i_c[701],c_t[701],s_t[701]);
fa fau_0_702(a_i_c[702],a_i_s[702],b_i_c[702],c_t[702],s_t[702]);
fa fau_0_703(a_i_c[703],a_i_s[703],b_i_c[703],c_t[703],s_t[703]);
fa fau_0_704(a_i_c[704],a_i_s[704],b_i_c[704],c_t[704],s_t[704]);
fa fau_0_705(a_i_c[705],a_i_s[705],b_i_c[705],c_t[705],s_t[705]);
fa fau_0_706(a_i_c[706],a_i_s[706],b_i_c[706],c_t[706],s_t[706]);
fa fau_0_707(a_i_c[707],a_i_s[707],b_i_c[707],c_t[707],s_t[707]);
fa fau_0_708(a_i_c[708],a_i_s[708],b_i_c[708],c_t[708],s_t[708]);
fa fau_0_709(a_i_c[709],a_i_s[709],b_i_c[709],c_t[709],s_t[709]);
fa fau_0_710(a_i_c[710],a_i_s[710],b_i_c[710],c_t[710],s_t[710]);
fa fau_0_711(a_i_c[711],a_i_s[711],b_i_c[711],c_t[711],s_t[711]);
fa fau_0_712(a_i_c[712],a_i_s[712],b_i_c[712],c_t[712],s_t[712]);
fa fau_0_713(a_i_c[713],a_i_s[713],b_i_c[713],c_t[713],s_t[713]);
fa fau_0_714(a_i_c[714],a_i_s[714],b_i_c[714],c_t[714],s_t[714]);
fa fau_0_715(a_i_c[715],a_i_s[715],b_i_c[715],c_t[715],s_t[715]);
fa fau_0_716(a_i_c[716],a_i_s[716],b_i_c[716],c_t[716],s_t[716]);
fa fau_0_717(a_i_c[717],a_i_s[717],b_i_c[717],c_t[717],s_t[717]);
fa fau_0_718(a_i_c[718],a_i_s[718],b_i_c[718],c_t[718],s_t[718]);
fa fau_0_719(a_i_c[719],a_i_s[719],b_i_c[719],c_t[719],s_t[719]);
fa fau_0_720(a_i_c[720],a_i_s[720],b_i_c[720],c_t[720],s_t[720]);
fa fau_0_721(a_i_c[721],a_i_s[721],b_i_c[721],c_t[721],s_t[721]);
fa fau_0_722(a_i_c[722],a_i_s[722],b_i_c[722],c_t[722],s_t[722]);
fa fau_0_723(a_i_c[723],a_i_s[723],b_i_c[723],c_t[723],s_t[723]);
fa fau_0_724(a_i_c[724],a_i_s[724],b_i_c[724],c_t[724],s_t[724]);
fa fau_0_725(a_i_c[725],a_i_s[725],b_i_c[725],c_t[725],s_t[725]);
fa fau_0_726(a_i_c[726],a_i_s[726],b_i_c[726],c_t[726],s_t[726]);
fa fau_0_727(a_i_c[727],a_i_s[727],b_i_c[727],c_t[727],s_t[727]);
fa fau_0_728(a_i_c[728],a_i_s[728],b_i_c[728],c_t[728],s_t[728]);
fa fau_0_729(a_i_c[729],a_i_s[729],b_i_c[729],c_t[729],s_t[729]);
fa fau_0_730(a_i_c[730],a_i_s[730],b_i_c[730],c_t[730],s_t[730]);
fa fau_0_731(a_i_c[731],a_i_s[731],b_i_c[731],c_t[731],s_t[731]);
fa fau_0_732(a_i_c[732],a_i_s[732],b_i_c[732],c_t[732],s_t[732]);
fa fau_0_733(a_i_c[733],a_i_s[733],b_i_c[733],c_t[733],s_t[733]);
fa fau_0_734(a_i_c[734],a_i_s[734],b_i_c[734],c_t[734],s_t[734]);
fa fau_0_735(a_i_c[735],a_i_s[735],b_i_c[735],c_t[735],s_t[735]);
fa fau_0_736(a_i_c[736],a_i_s[736],b_i_c[736],c_t[736],s_t[736]);
fa fau_0_737(a_i_c[737],a_i_s[737],b_i_c[737],c_t[737],s_t[737]);
fa fau_0_738(a_i_c[738],a_i_s[738],b_i_c[738],c_t[738],s_t[738]);
fa fau_0_739(a_i_c[739],a_i_s[739],b_i_c[739],c_t[739],s_t[739]);
fa fau_0_740(a_i_c[740],a_i_s[740],b_i_c[740],c_t[740],s_t[740]);
fa fau_0_741(a_i_c[741],a_i_s[741],b_i_c[741],c_t[741],s_t[741]);
fa fau_0_742(a_i_c[742],a_i_s[742],b_i_c[742],c_t[742],s_t[742]);
fa fau_0_743(a_i_c[743],a_i_s[743],b_i_c[743],c_t[743],s_t[743]);
fa fau_0_744(a_i_c[744],a_i_s[744],b_i_c[744],c_t[744],s_t[744]);
fa fau_0_745(a_i_c[745],a_i_s[745],b_i_c[745],c_t[745],s_t[745]);
fa fau_0_746(a_i_c[746],a_i_s[746],b_i_c[746],c_t[746],s_t[746]);
fa fau_0_747(a_i_c[747],a_i_s[747],b_i_c[747],c_t[747],s_t[747]);
fa fau_0_748(a_i_c[748],a_i_s[748],b_i_c[748],c_t[748],s_t[748]);
fa fau_0_749(a_i_c[749],a_i_s[749],b_i_c[749],c_t[749],s_t[749]);
fa fau_0_750(a_i_c[750],a_i_s[750],b_i_c[750],c_t[750],s_t[750]);
fa fau_0_751(a_i_c[751],a_i_s[751],b_i_c[751],c_t[751],s_t[751]);
fa fau_0_752(a_i_c[752],a_i_s[752],b_i_c[752],c_t[752],s_t[752]);
fa fau_0_753(a_i_c[753],a_i_s[753],b_i_c[753],c_t[753],s_t[753]);
fa fau_0_754(a_i_c[754],a_i_s[754],b_i_c[754],c_t[754],s_t[754]);
fa fau_0_755(a_i_c[755],a_i_s[755],b_i_c[755],c_t[755],s_t[755]);
fa fau_0_756(a_i_c[756],a_i_s[756],b_i_c[756],c_t[756],s_t[756]);
fa fau_0_757(a_i_c[757],a_i_s[757],b_i_c[757],c_t[757],s_t[757]);
fa fau_0_758(a_i_c[758],a_i_s[758],b_i_c[758],c_t[758],s_t[758]);
fa fau_0_759(a_i_c[759],a_i_s[759],b_i_c[759],c_t[759],s_t[759]);
fa fau_0_760(a_i_c[760],a_i_s[760],b_i_c[760],c_t[760],s_t[760]);
fa fau_0_761(a_i_c[761],a_i_s[761],b_i_c[761],c_t[761],s_t[761]);
fa fau_0_762(a_i_c[762],a_i_s[762],b_i_c[762],c_t[762],s_t[762]);
fa fau_0_763(a_i_c[763],a_i_s[763],b_i_c[763],c_t[763],s_t[763]);
fa fau_0_764(a_i_c[764],a_i_s[764],b_i_c[764],c_t[764],s_t[764]);
fa fau_0_765(a_i_c[765],a_i_s[765],b_i_c[765],c_t[765],s_t[765]);
fa fau_0_766(a_i_c[766],a_i_s[766],b_i_c[766],c_t[766],s_t[766]);
fa fau_0_767(a_i_c[767],a_i_s[767],b_i_c[767],c_t[767],s_t[767]);
fa fau_0_768(a_i_c[768],a_i_s[768],b_i_c[768],c_t[768],s_t[768]);
fa fau_0_769(a_i_c[769],a_i_s[769],b_i_c[769],c_t[769],s_t[769]);
fa fau_0_770(a_i_c[770],a_i_s[770],b_i_c[770],c_t[770],s_t[770]);
fa fau_0_771(a_i_c[771],a_i_s[771],b_i_c[771],c_t[771],s_t[771]);
fa fau_0_772(a_i_c[772],a_i_s[772],b_i_c[772],c_t[772],s_t[772]);
fa fau_0_773(a_i_c[773],a_i_s[773],b_i_c[773],c_t[773],s_t[773]);
fa fau_0_774(a_i_c[774],a_i_s[774],b_i_c[774],c_t[774],s_t[774]);
fa fau_0_775(a_i_c[775],a_i_s[775],b_i_c[775],c_t[775],s_t[775]);
fa fau_0_776(a_i_c[776],a_i_s[776],b_i_c[776],c_t[776],s_t[776]);
fa fau_0_777(a_i_c[777],a_i_s[777],b_i_c[777],c_t[777],s_t[777]);
fa fau_0_778(a_i_c[778],a_i_s[778],b_i_c[778],c_t[778],s_t[778]);
fa fau_0_779(a_i_c[779],a_i_s[779],b_i_c[779],c_t[779],s_t[779]);
fa fau_0_780(a_i_c[780],a_i_s[780],b_i_c[780],c_t[780],s_t[780]);
fa fau_0_781(a_i_c[781],a_i_s[781],b_i_c[781],c_t[781],s_t[781]);
fa fau_0_782(a_i_c[782],a_i_s[782],b_i_c[782],c_t[782],s_t[782]);
fa fau_0_783(a_i_c[783],a_i_s[783],b_i_c[783],c_t[783],s_t[783]);
fa fau_0_784(a_i_c[784],a_i_s[784],b_i_c[784],c_t[784],s_t[784]);
fa fau_0_785(a_i_c[785],a_i_s[785],b_i_c[785],c_t[785],s_t[785]);
fa fau_0_786(a_i_c[786],a_i_s[786],b_i_c[786],c_t[786],s_t[786]);
fa fau_0_787(a_i_c[787],a_i_s[787],b_i_c[787],c_t[787],s_t[787]);
fa fau_0_788(a_i_c[788],a_i_s[788],b_i_c[788],c_t[788],s_t[788]);
fa fau_0_789(a_i_c[789],a_i_s[789],b_i_c[789],c_t[789],s_t[789]);
fa fau_0_790(a_i_c[790],a_i_s[790],b_i_c[790],c_t[790],s_t[790]);
fa fau_0_791(a_i_c[791],a_i_s[791],b_i_c[791],c_t[791],s_t[791]);
fa fau_0_792(a_i_c[792],a_i_s[792],b_i_c[792],c_t[792],s_t[792]);
fa fau_0_793(a_i_c[793],a_i_s[793],b_i_c[793],c_t[793],s_t[793]);
fa fau_0_794(a_i_c[794],a_i_s[794],b_i_c[794],c_t[794],s_t[794]);
fa fau_0_795(a_i_c[795],a_i_s[795],b_i_c[795],c_t[795],s_t[795]);
fa fau_0_796(a_i_c[796],a_i_s[796],b_i_c[796],c_t[796],s_t[796]);
fa fau_0_797(a_i_c[797],a_i_s[797],b_i_c[797],c_t[797],s_t[797]);
fa fau_0_798(a_i_c[798],a_i_s[798],b_i_c[798],c_t[798],s_t[798]);
fa fau_0_799(a_i_c[799],a_i_s[799],b_i_c[799],c_t[799],s_t[799]);
fa fau_0_800(a_i_c[800],a_i_s[800],b_i_c[800],c_t[800],s_t[800]);
fa fau_0_801(a_i_c[801],a_i_s[801],b_i_c[801],c_t[801],s_t[801]);
fa fau_0_802(a_i_c[802],a_i_s[802],b_i_c[802],c_t[802],s_t[802]);
fa fau_0_803(a_i_c[803],a_i_s[803],b_i_c[803],c_t[803],s_t[803]);
fa fau_0_804(a_i_c[804],a_i_s[804],b_i_c[804],c_t[804],s_t[804]);
fa fau_0_805(a_i_c[805],a_i_s[805],b_i_c[805],c_t[805],s_t[805]);
fa fau_0_806(a_i_c[806],a_i_s[806],b_i_c[806],c_t[806],s_t[806]);
fa fau_0_807(a_i_c[807],a_i_s[807],b_i_c[807],c_t[807],s_t[807]);
fa fau_0_808(a_i_c[808],a_i_s[808],b_i_c[808],c_t[808],s_t[808]);
fa fau_0_809(a_i_c[809],a_i_s[809],b_i_c[809],c_t[809],s_t[809]);
fa fau_0_810(a_i_c[810],a_i_s[810],b_i_c[810],c_t[810],s_t[810]);
fa fau_0_811(a_i_c[811],a_i_s[811],b_i_c[811],c_t[811],s_t[811]);
fa fau_0_812(a_i_c[812],a_i_s[812],b_i_c[812],c_t[812],s_t[812]);
fa fau_0_813(a_i_c[813],a_i_s[813],b_i_c[813],c_t[813],s_t[813]);
fa fau_0_814(a_i_c[814],a_i_s[814],b_i_c[814],c_t[814],s_t[814]);
fa fau_0_815(a_i_c[815],a_i_s[815],b_i_c[815],c_t[815],s_t[815]);
fa fau_0_816(a_i_c[816],a_i_s[816],b_i_c[816],c_t[816],s_t[816]);
fa fau_0_817(a_i_c[817],a_i_s[817],b_i_c[817],c_t[817],s_t[817]);
fa fau_0_818(a_i_c[818],a_i_s[818],b_i_c[818],c_t[818],s_t[818]);
fa fau_0_819(a_i_c[819],a_i_s[819],b_i_c[819],c_t[819],s_t[819]);
fa fau_0_820(a_i_c[820],a_i_s[820],b_i_c[820],c_t[820],s_t[820]);
fa fau_0_821(a_i_c[821],a_i_s[821],b_i_c[821],c_t[821],s_t[821]);
fa fau_0_822(a_i_c[822],a_i_s[822],b_i_c[822],c_t[822],s_t[822]);
fa fau_0_823(a_i_c[823],a_i_s[823],b_i_c[823],c_t[823],s_t[823]);
fa fau_0_824(a_i_c[824],a_i_s[824],b_i_c[824],c_t[824],s_t[824]);
fa fau_0_825(a_i_c[825],a_i_s[825],b_i_c[825],c_t[825],s_t[825]);
fa fau_0_826(a_i_c[826],a_i_s[826],b_i_c[826],c_t[826],s_t[826]);
fa fau_0_827(a_i_c[827],a_i_s[827],b_i_c[827],c_t[827],s_t[827]);
fa fau_0_828(a_i_c[828],a_i_s[828],b_i_c[828],c_t[828],s_t[828]);
fa fau_0_829(a_i_c[829],a_i_s[829],b_i_c[829],c_t[829],s_t[829]);
fa fau_0_830(a_i_c[830],a_i_s[830],b_i_c[830],c_t[830],s_t[830]);
fa fau_0_831(a_i_c[831],a_i_s[831],b_i_c[831],c_t[831],s_t[831]);
fa fau_0_832(a_i_c[832],a_i_s[832],b_i_c[832],c_t[832],s_t[832]);
fa fau_0_833(a_i_c[833],a_i_s[833],b_i_c[833],c_t[833],s_t[833]);
fa fau_0_834(a_i_c[834],a_i_s[834],b_i_c[834],c_t[834],s_t[834]);
fa fau_0_835(a_i_c[835],a_i_s[835],b_i_c[835],c_t[835],s_t[835]);
fa fau_0_836(a_i_c[836],a_i_s[836],b_i_c[836],c_t[836],s_t[836]);
fa fau_0_837(a_i_c[837],a_i_s[837],b_i_c[837],c_t[837],s_t[837]);
fa fau_0_838(a_i_c[838],a_i_s[838],b_i_c[838],c_t[838],s_t[838]);
fa fau_0_839(a_i_c[839],a_i_s[839],b_i_c[839],c_t[839],s_t[839]);
fa fau_0_840(a_i_c[840],a_i_s[840],b_i_c[840],c_t[840],s_t[840]);
fa fau_0_841(a_i_c[841],a_i_s[841],b_i_c[841],c_t[841],s_t[841]);
fa fau_0_842(a_i_c[842],a_i_s[842],b_i_c[842],c_t[842],s_t[842]);
fa fau_0_843(a_i_c[843],a_i_s[843],b_i_c[843],c_t[843],s_t[843]);
fa fau_0_844(a_i_c[844],a_i_s[844],b_i_c[844],c_t[844],s_t[844]);
fa fau_0_845(a_i_c[845],a_i_s[845],b_i_c[845],c_t[845],s_t[845]);
fa fau_0_846(a_i_c[846],a_i_s[846],b_i_c[846],c_t[846],s_t[846]);
fa fau_0_847(a_i_c[847],a_i_s[847],b_i_c[847],c_t[847],s_t[847]);
fa fau_0_848(a_i_c[848],a_i_s[848],b_i_c[848],c_t[848],s_t[848]);
fa fau_0_849(a_i_c[849],a_i_s[849],b_i_c[849],c_t[849],s_t[849]);
fa fau_0_850(a_i_c[850],a_i_s[850],b_i_c[850],c_t[850],s_t[850]);
fa fau_0_851(a_i_c[851],a_i_s[851],b_i_c[851],c_t[851],s_t[851]);
fa fau_0_852(a_i_c[852],a_i_s[852],b_i_c[852],c_t[852],s_t[852]);
fa fau_0_853(a_i_c[853],a_i_s[853],b_i_c[853],c_t[853],s_t[853]);
fa fau_0_854(a_i_c[854],a_i_s[854],b_i_c[854],c_t[854],s_t[854]);
fa fau_0_855(a_i_c[855],a_i_s[855],b_i_c[855],c_t[855],s_t[855]);
fa fau_0_856(a_i_c[856],a_i_s[856],b_i_c[856],c_t[856],s_t[856]);
fa fau_0_857(a_i_c[857],a_i_s[857],b_i_c[857],c_t[857],s_t[857]);
fa fau_0_858(a_i_c[858],a_i_s[858],b_i_c[858],c_t[858],s_t[858]);
fa fau_0_859(a_i_c[859],a_i_s[859],b_i_c[859],c_t[859],s_t[859]);
fa fau_0_860(a_i_c[860],a_i_s[860],b_i_c[860],c_t[860],s_t[860]);
fa fau_0_861(a_i_c[861],a_i_s[861],b_i_c[861],c_t[861],s_t[861]);
fa fau_0_862(a_i_c[862],a_i_s[862],b_i_c[862],c_t[862],s_t[862]);
fa fau_0_863(a_i_c[863],a_i_s[863],b_i_c[863],c_t[863],s_t[863]);
fa fau_0_864(a_i_c[864],a_i_s[864],b_i_c[864],c_t[864],s_t[864]);
fa fau_0_865(a_i_c[865],a_i_s[865],b_i_c[865],c_t[865],s_t[865]);
fa fau_0_866(a_i_c[866],a_i_s[866],b_i_c[866],c_t[866],s_t[866]);
fa fau_0_867(a_i_c[867],a_i_s[867],b_i_c[867],c_t[867],s_t[867]);
fa fau_0_868(a_i_c[868],a_i_s[868],b_i_c[868],c_t[868],s_t[868]);
fa fau_0_869(a_i_c[869],a_i_s[869],b_i_c[869],c_t[869],s_t[869]);
fa fau_0_870(a_i_c[870],a_i_s[870],b_i_c[870],c_t[870],s_t[870]);
fa fau_0_871(a_i_c[871],a_i_s[871],b_i_c[871],c_t[871],s_t[871]);
fa fau_0_872(a_i_c[872],a_i_s[872],b_i_c[872],c_t[872],s_t[872]);
fa fau_0_873(a_i_c[873],a_i_s[873],b_i_c[873],c_t[873],s_t[873]);
fa fau_0_874(a_i_c[874],a_i_s[874],b_i_c[874],c_t[874],s_t[874]);
fa fau_0_875(a_i_c[875],a_i_s[875],b_i_c[875],c_t[875],s_t[875]);
fa fau_0_876(a_i_c[876],a_i_s[876],b_i_c[876],c_t[876],s_t[876]);
fa fau_0_877(a_i_c[877],a_i_s[877],b_i_c[877],c_t[877],s_t[877]);
fa fau_0_878(a_i_c[878],a_i_s[878],b_i_c[878],c_t[878],s_t[878]);
fa fau_0_879(a_i_c[879],a_i_s[879],b_i_c[879],c_t[879],s_t[879]);
fa fau_0_880(a_i_c[880],a_i_s[880],b_i_c[880],c_t[880],s_t[880]);
fa fau_0_881(a_i_c[881],a_i_s[881],b_i_c[881],c_t[881],s_t[881]);
fa fau_0_882(a_i_c[882],a_i_s[882],b_i_c[882],c_t[882],s_t[882]);
fa fau_0_883(a_i_c[883],a_i_s[883],b_i_c[883],c_t[883],s_t[883]);
fa fau_0_884(a_i_c[884],a_i_s[884],b_i_c[884],c_t[884],s_t[884]);
fa fau_0_885(a_i_c[885],a_i_s[885],b_i_c[885],c_t[885],s_t[885]);
fa fau_0_886(a_i_c[886],a_i_s[886],b_i_c[886],c_t[886],s_t[886]);
fa fau_0_887(a_i_c[887],a_i_s[887],b_i_c[887],c_t[887],s_t[887]);
fa fau_0_888(a_i_c[888],a_i_s[888],b_i_c[888],c_t[888],s_t[888]);
fa fau_0_889(a_i_c[889],a_i_s[889],b_i_c[889],c_t[889],s_t[889]);
fa fau_0_890(a_i_c[890],a_i_s[890],b_i_c[890],c_t[890],s_t[890]);
fa fau_0_891(a_i_c[891],a_i_s[891],b_i_c[891],c_t[891],s_t[891]);
fa fau_0_892(a_i_c[892],a_i_s[892],b_i_c[892],c_t[892],s_t[892]);
fa fau_0_893(a_i_c[893],a_i_s[893],b_i_c[893],c_t[893],s_t[893]);
fa fau_0_894(a_i_c[894],a_i_s[894],b_i_c[894],c_t[894],s_t[894]);
fa fau_0_895(a_i_c[895],a_i_s[895],b_i_c[895],c_t[895],s_t[895]);
fa fau_0_896(a_i_c[896],a_i_s[896],b_i_c[896],c_t[896],s_t[896]);
fa fau_0_897(a_i_c[897],a_i_s[897],b_i_c[897],c_t[897],s_t[897]);
fa fau_0_898(a_i_c[898],a_i_s[898],b_i_c[898],c_t[898],s_t[898]);
fa fau_0_899(a_i_c[899],a_i_s[899],b_i_c[899],c_t[899],s_t[899]);
fa fau_0_900(a_i_c[900],a_i_s[900],b_i_c[900],c_t[900],s_t[900]);
fa fau_0_901(a_i_c[901],a_i_s[901],b_i_c[901],c_t[901],s_t[901]);
fa fau_0_902(a_i_c[902],a_i_s[902],b_i_c[902],c_t[902],s_t[902]);
fa fau_0_903(a_i_c[903],a_i_s[903],b_i_c[903],c_t[903],s_t[903]);
fa fau_0_904(a_i_c[904],a_i_s[904],b_i_c[904],c_t[904],s_t[904]);
fa fau_0_905(a_i_c[905],a_i_s[905],b_i_c[905],c_t[905],s_t[905]);
fa fau_0_906(a_i_c[906],a_i_s[906],b_i_c[906],c_t[906],s_t[906]);
fa fau_0_907(a_i_c[907],a_i_s[907],b_i_c[907],c_t[907],s_t[907]);
fa fau_0_908(a_i_c[908],a_i_s[908],b_i_c[908],c_t[908],s_t[908]);
fa fau_0_909(a_i_c[909],a_i_s[909],b_i_c[909],c_t[909],s_t[909]);
fa fau_0_910(a_i_c[910],a_i_s[910],b_i_c[910],c_t[910],s_t[910]);
fa fau_0_911(a_i_c[911],a_i_s[911],b_i_c[911],c_t[911],s_t[911]);
fa fau_0_912(a_i_c[912],a_i_s[912],b_i_c[912],c_t[912],s_t[912]);
fa fau_0_913(a_i_c[913],a_i_s[913],b_i_c[913],c_t[913],s_t[913]);
fa fau_0_914(a_i_c[914],a_i_s[914],b_i_c[914],c_t[914],s_t[914]);
fa fau_0_915(a_i_c[915],a_i_s[915],b_i_c[915],c_t[915],s_t[915]);
fa fau_0_916(a_i_c[916],a_i_s[916],b_i_c[916],c_t[916],s_t[916]);
fa fau_0_917(a_i_c[917],a_i_s[917],b_i_c[917],c_t[917],s_t[917]);
fa fau_0_918(a_i_c[918],a_i_s[918],b_i_c[918],c_t[918],s_t[918]);
fa fau_0_919(a_i_c[919],a_i_s[919],b_i_c[919],c_t[919],s_t[919]);
fa fau_0_920(a_i_c[920],a_i_s[920],b_i_c[920],c_t[920],s_t[920]);
fa fau_0_921(a_i_c[921],a_i_s[921],b_i_c[921],c_t[921],s_t[921]);
fa fau_0_922(a_i_c[922],a_i_s[922],b_i_c[922],c_t[922],s_t[922]);
fa fau_0_923(a_i_c[923],a_i_s[923],b_i_c[923],c_t[923],s_t[923]);
fa fau_0_924(a_i_c[924],a_i_s[924],b_i_c[924],c_t[924],s_t[924]);
fa fau_0_925(a_i_c[925],a_i_s[925],b_i_c[925],c_t[925],s_t[925]);
fa fau_0_926(a_i_c[926],a_i_s[926],b_i_c[926],c_t[926],s_t[926]);
fa fau_0_927(a_i_c[927],a_i_s[927],b_i_c[927],c_t[927],s_t[927]);
fa fau_0_928(a_i_c[928],a_i_s[928],b_i_c[928],c_t[928],s_t[928]);
fa fau_0_929(a_i_c[929],a_i_s[929],b_i_c[929],c_t[929],s_t[929]);
fa fau_0_930(a_i_c[930],a_i_s[930],b_i_c[930],c_t[930],s_t[930]);
fa fau_0_931(a_i_c[931],a_i_s[931],b_i_c[931],c_t[931],s_t[931]);
fa fau_0_932(a_i_c[932],a_i_s[932],b_i_c[932],c_t[932],s_t[932]);
fa fau_0_933(a_i_c[933],a_i_s[933],b_i_c[933],c_t[933],s_t[933]);
fa fau_0_934(a_i_c[934],a_i_s[934],b_i_c[934],c_t[934],s_t[934]);
fa fau_0_935(a_i_c[935],a_i_s[935],b_i_c[935],c_t[935],s_t[935]);
fa fau_0_936(a_i_c[936],a_i_s[936],b_i_c[936],c_t[936],s_t[936]);
fa fau_0_937(a_i_c[937],a_i_s[937],b_i_c[937],c_t[937],s_t[937]);
fa fau_0_938(a_i_c[938],a_i_s[938],b_i_c[938],c_t[938],s_t[938]);
fa fau_0_939(a_i_c[939],a_i_s[939],b_i_c[939],c_t[939],s_t[939]);
fa fau_0_940(a_i_c[940],a_i_s[940],b_i_c[940],c_t[940],s_t[940]);
fa fau_0_941(a_i_c[941],a_i_s[941],b_i_c[941],c_t[941],s_t[941]);
fa fau_0_942(a_i_c[942],a_i_s[942],b_i_c[942],c_t[942],s_t[942]);
fa fau_0_943(a_i_c[943],a_i_s[943],b_i_c[943],c_t[943],s_t[943]);
fa fau_0_944(a_i_c[944],a_i_s[944],b_i_c[944],c_t[944],s_t[944]);
fa fau_0_945(a_i_c[945],a_i_s[945],b_i_c[945],c_t[945],s_t[945]);
fa fau_0_946(a_i_c[946],a_i_s[946],b_i_c[946],c_t[946],s_t[946]);
fa fau_0_947(a_i_c[947],a_i_s[947],b_i_c[947],c_t[947],s_t[947]);
fa fau_0_948(a_i_c[948],a_i_s[948],b_i_c[948],c_t[948],s_t[948]);
fa fau_0_949(a_i_c[949],a_i_s[949],b_i_c[949],c_t[949],s_t[949]);
fa fau_0_950(a_i_c[950],a_i_s[950],b_i_c[950],c_t[950],s_t[950]);
fa fau_0_951(a_i_c[951],a_i_s[951],b_i_c[951],c_t[951],s_t[951]);
fa fau_0_952(a_i_c[952],a_i_s[952],b_i_c[952],c_t[952],s_t[952]);
fa fau_0_953(a_i_c[953],a_i_s[953],b_i_c[953],c_t[953],s_t[953]);
fa fau_0_954(a_i_c[954],a_i_s[954],b_i_c[954],c_t[954],s_t[954]);
fa fau_0_955(a_i_c[955],a_i_s[955],b_i_c[955],c_t[955],s_t[955]);
fa fau_0_956(a_i_c[956],a_i_s[956],b_i_c[956],c_t[956],s_t[956]);
fa fau_0_957(a_i_c[957],a_i_s[957],b_i_c[957],c_t[957],s_t[957]);
fa fau_0_958(a_i_c[958],a_i_s[958],b_i_c[958],c_t[958],s_t[958]);
fa fau_0_959(a_i_c[959],a_i_s[959],b_i_c[959],c_t[959],s_t[959]);
fa fau_0_960(a_i_c[960],a_i_s[960],b_i_c[960],c_t[960],s_t[960]);
fa fau_0_961(a_i_c[961],a_i_s[961],b_i_c[961],c_t[961],s_t[961]);
fa fau_0_962(a_i_c[962],a_i_s[962],b_i_c[962],c_t[962],s_t[962]);
fa fau_0_963(a_i_c[963],a_i_s[963],b_i_c[963],c_t[963],s_t[963]);
fa fau_0_964(a_i_c[964],a_i_s[964],b_i_c[964],c_t[964],s_t[964]);
fa fau_0_965(a_i_c[965],a_i_s[965],b_i_c[965],c_t[965],s_t[965]);
fa fau_0_966(a_i_c[966],a_i_s[966],b_i_c[966],c_t[966],s_t[966]);
fa fau_0_967(a_i_c[967],a_i_s[967],b_i_c[967],c_t[967],s_t[967]);
fa fau_0_968(a_i_c[968],a_i_s[968],b_i_c[968],c_t[968],s_t[968]);
fa fau_0_969(a_i_c[969],a_i_s[969],b_i_c[969],c_t[969],s_t[969]);
fa fau_0_970(a_i_c[970],a_i_s[970],b_i_c[970],c_t[970],s_t[970]);
fa fau_0_971(a_i_c[971],a_i_s[971],b_i_c[971],c_t[971],s_t[971]);
fa fau_0_972(a_i_c[972],a_i_s[972],b_i_c[972],c_t[972],s_t[972]);
fa fau_0_973(a_i_c[973],a_i_s[973],b_i_c[973],c_t[973],s_t[973]);
fa fau_0_974(a_i_c[974],a_i_s[974],b_i_c[974],c_t[974],s_t[974]);
fa fau_0_975(a_i_c[975],a_i_s[975],b_i_c[975],c_t[975],s_t[975]);
fa fau_0_976(a_i_c[976],a_i_s[976],b_i_c[976],c_t[976],s_t[976]);
fa fau_0_977(a_i_c[977],a_i_s[977],b_i_c[977],c_t[977],s_t[977]);
fa fau_0_978(a_i_c[978],a_i_s[978],b_i_c[978],c_t[978],s_t[978]);
fa fau_0_979(a_i_c[979],a_i_s[979],b_i_c[979],c_t[979],s_t[979]);
fa fau_0_980(a_i_c[980],a_i_s[980],b_i_c[980],c_t[980],s_t[980]);
fa fau_0_981(a_i_c[981],a_i_s[981],b_i_c[981],c_t[981],s_t[981]);
fa fau_0_982(a_i_c[982],a_i_s[982],b_i_c[982],c_t[982],s_t[982]);
fa fau_0_983(a_i_c[983],a_i_s[983],b_i_c[983],c_t[983],s_t[983]);
fa fau_0_984(a_i_c[984],a_i_s[984],b_i_c[984],c_t[984],s_t[984]);
fa fau_0_985(a_i_c[985],a_i_s[985],b_i_c[985],c_t[985],s_t[985]);
fa fau_0_986(a_i_c[986],a_i_s[986],b_i_c[986],c_t[986],s_t[986]);
fa fau_0_987(a_i_c[987],a_i_s[987],b_i_c[987],c_t[987],s_t[987]);
fa fau_0_988(a_i_c[988],a_i_s[988],b_i_c[988],c_t[988],s_t[988]);
fa fau_0_989(a_i_c[989],a_i_s[989],b_i_c[989],c_t[989],s_t[989]);
fa fau_0_990(a_i_c[990],a_i_s[990],b_i_c[990],c_t[990],s_t[990]);
fa fau_0_991(a_i_c[991],a_i_s[991],b_i_c[991],c_t[991],s_t[991]);
fa fau_0_992(a_i_c[992],a_i_s[992],b_i_c[992],c_t[992],s_t[992]);
fa fau_0_993(a_i_c[993],a_i_s[993],b_i_c[993],c_t[993],s_t[993]);
fa fau_0_994(a_i_c[994],a_i_s[994],b_i_c[994],c_t[994],s_t[994]);
fa fau_0_995(a_i_c[995],a_i_s[995],b_i_c[995],c_t[995],s_t[995]);
fa fau_0_996(a_i_c[996],a_i_s[996],b_i_c[996],c_t[996],s_t[996]);
fa fau_0_997(a_i_c[997],a_i_s[997],b_i_c[997],c_t[997],s_t[997]);
fa fau_0_998(a_i_c[998],a_i_s[998],b_i_c[998],c_t[998],s_t[998]);
fa fau_0_999(a_i_c[999],a_i_s[999],b_i_c[999],c_t[999],s_t[999]);
fa fau_0_1000(a_i_c[1000],a_i_s[1000],b_i_c[1000],c_t[1000],s_t[1000]);
fa fau_0_1001(a_i_c[1001],a_i_s[1001],b_i_c[1001],c_t[1001],s_t[1001]);
fa fau_0_1002(a_i_c[1002],a_i_s[1002],b_i_c[1002],c_t[1002],s_t[1002]);
fa fau_0_1003(a_i_c[1003],a_i_s[1003],b_i_c[1003],c_t[1003],s_t[1003]);
fa fau_0_1004(a_i_c[1004],a_i_s[1004],b_i_c[1004],c_t[1004],s_t[1004]);
fa fau_0_1005(a_i_c[1005],a_i_s[1005],b_i_c[1005],c_t[1005],s_t[1005]);
fa fau_0_1006(a_i_c[1006],a_i_s[1006],b_i_c[1006],c_t[1006],s_t[1006]);
fa fau_0_1007(a_i_c[1007],a_i_s[1007],b_i_c[1007],c_t[1007],s_t[1007]);
fa fau_0_1008(a_i_c[1008],a_i_s[1008],b_i_c[1008],c_t[1008],s_t[1008]);
fa fau_0_1009(a_i_c[1009],a_i_s[1009],b_i_c[1009],c_t[1009],s_t[1009]);
fa fau_0_1010(a_i_c[1010],a_i_s[1010],b_i_c[1010],c_t[1010],s_t[1010]);
fa fau_0_1011(a_i_c[1011],a_i_s[1011],b_i_c[1011],c_t[1011],s_t[1011]);
fa fau_0_1012(a_i_c[1012],a_i_s[1012],b_i_c[1012],c_t[1012],s_t[1012]);
fa fau_0_1013(a_i_c[1013],a_i_s[1013],b_i_c[1013],c_t[1013],s_t[1013]);
fa fau_0_1014(a_i_c[1014],a_i_s[1014],b_i_c[1014],c_t[1014],s_t[1014]);
fa fau_0_1015(a_i_c[1015],a_i_s[1015],b_i_c[1015],c_t[1015],s_t[1015]);
fa fau_0_1016(a_i_c[1016],a_i_s[1016],b_i_c[1016],c_t[1016],s_t[1016]);
fa fau_0_1017(a_i_c[1017],a_i_s[1017],b_i_c[1017],c_t[1017],s_t[1017]);
fa fau_0_1018(a_i_c[1018],a_i_s[1018],b_i_c[1018],c_t[1018],s_t[1018]);
fa fau_0_1019(a_i_c[1019],a_i_s[1019],b_i_c[1019],c_t[1019],s_t[1019]);
fa fau_0_1020(a_i_c[1020],a_i_s[1020],b_i_c[1020],c_t[1020],s_t[1020]);
fa fau_0_1021(a_i_c[1021],a_i_s[1021],b_i_c[1021],c_t[1021],s_t[1021]);
fa fau_0_1022(a_i_c[1022],a_i_s[1022],b_i_c[1022],c_t[1022],s_t[1022]);
fa fau_0_1023(a_i_c[1023],a_i_s[1023],b_i_c[1023],c_t[1023],s_t[1023]);
fa fau_0_1024(a_i_c[1024],a_i_s[1024],b_i_c[1024],c_t[1024],s_t[1024]);
fa fau_0_1025(a_i_c[1025],a_i_s[1025],b_i_c[1025],c_t[1025],s_t[1025]);
fa fau_0_1026(a_i_c[1026],a_i_s[1026],b_i_c[1026],c_t[1026],s_t[1026]);
fa fau_0_1027(a_i_c[1027],a_i_s[1027],b_i_c[1027],c_t[1027],s_t[1027]);
fa fau_0_1028(a_i_c[1028],a_i_s[1028],b_i_c[1028],c_t[1028],s_t[1028]);
fa fau_0_1029(a_i_c[1029],a_i_s[1029],b_i_c[1029],c_t[1029],s_t[1029]);
fa fau_0_1030(a_i_c[1030],a_i_s[1030],b_i_c[1030],c_t[1030],s_t[1030]);
fa fau_0_1031(a_i_c[1031],a_i_s[1031],b_i_c[1031],c_t[1031],s_t[1031]);
fa fau_0_1032(a_i_c[1032],a_i_s[1032],b_i_c[1032],c_t[1032],s_t[1032]);
fa fau_0_1033(a_i_c[1033],a_i_s[1033],b_i_c[1033],c_t[1033],s_t[1033]);
fa fau_0_1034(a_i_c[1034],a_i_s[1034],b_i_c[1034],c_t[1034],s_t[1034]);
fa fau_0_1035(a_i_c[1035],a_i_s[1035],b_i_c[1035],c_t[1035],s_t[1035]);
fa fau_0_1036(a_i_c[1036],a_i_s[1036],b_i_c[1036],c_t[1036],s_t[1036]);
fa fau_0_1037(a_i_c[1037],a_i_s[1037],b_i_c[1037],c_t[1037],s_t[1037]);
fa fau_0_1038(a_i_c[1038],a_i_s[1038],b_i_c[1038],c_t[1038],s_t[1038]);
fa fau_0_1039(a_i_c[1039],a_i_s[1039],b_i_c[1039],c_t[1039],s_t[1039]);
fa fau_0_1040(a_i_c[1040],a_i_s[1040],b_i_c[1040],c_t[1040],s_t[1040]);
fa fau_0_1041(a_i_c[1041],a_i_s[1041],b_i_c[1041],c_t[1041],s_t[1041]);
fa fau_0_1042(a_i_c[1042],a_i_s[1042],b_i_c[1042],c_t[1042],s_t[1042]);
fa fau_0_1043(a_i_c[1043],a_i_s[1043],b_i_c[1043],c_t[1043],s_t[1043]);
fa fau_0_1044(a_i_c[1044],a_i_s[1044],b_i_c[1044],c_t[1044],s_t[1044]);
fa fau_0_1045(a_i_c[1045],a_i_s[1045],b_i_c[1045],c_t[1045],s_t[1045]);
fa fau_0_1046(a_i_c[1046],a_i_s[1046],b_i_c[1046],c_t[1046],s_t[1046]);
fa fau_0_1047(a_i_c[1047],a_i_s[1047],b_i_c[1047],c_t[1047],s_t[1047]);
fa fau_0_1048(a_i_c[1048],a_i_s[1048],b_i_c[1048],c_t[1048],s_t[1048]);
fa fau_0_1049(a_i_c[1049],a_i_s[1049],b_i_c[1049],c_t[1049],s_t[1049]);
fa fau_0_1050(a_i_c[1050],a_i_s[1050],b_i_c[1050],c_t[1050],s_t[1050]);
fa fau_0_1051(a_i_c[1051],a_i_s[1051],b_i_c[1051],c_t[1051],s_t[1051]);
fa fau_0_1052(a_i_c[1052],a_i_s[1052],b_i_c[1052],c_t[1052],s_t[1052]);
fa fau_0_1053(a_i_c[1053],a_i_s[1053],b_i_c[1053],c_t[1053],s_t[1053]);
fa fau_0_1054(a_i_c[1054],a_i_s[1054],b_i_c[1054],c_t[1054],s_t[1054]);
fa fau_0_1055(a_i_c[1055],a_i_s[1055],b_i_c[1055],c_t[1055],s_t[1055]);
fa fau_0_1056(a_i_c[1056],a_i_s[1056],b_i_c[1056],c_t[1056],s_t[1056]);
fa fau_0_1057(a_i_c[1057],a_i_s[1057],b_i_c[1057],c_t[1057],s_t[1057]);
fa fau_0_1058(a_i_c[1058],a_i_s[1058],b_i_c[1058],c_t[1058],s_t[1058]);
fa fau_0_1059(a_i_c[1059],a_i_s[1059],b_i_c[1059],c_t[1059],s_t[1059]);
fa fau_0_1060(a_i_c[1060],a_i_s[1060],b_i_c[1060],c_t[1060],s_t[1060]);
fa fau_0_1061(a_i_c[1061],a_i_s[1061],b_i_c[1061],c_t[1061],s_t[1061]);
fa fau_0_1062(a_i_c[1062],a_i_s[1062],b_i_c[1062],c_t[1062],s_t[1062]);
fa fau_0_1063(a_i_c[1063],a_i_s[1063],b_i_c[1063],c_t[1063],s_t[1063]);
fa fau_0_1064(a_i_c[1064],a_i_s[1064],b_i_c[1064],c_t[1064],s_t[1064]);
fa fau_0_1065(a_i_c[1065],a_i_s[1065],b_i_c[1065],c_t[1065],s_t[1065]);
fa fau_0_1066(a_i_c[1066],a_i_s[1066],b_i_c[1066],c_t[1066],s_t[1066]);
fa fau_0_1067(a_i_c[1067],a_i_s[1067],b_i_c[1067],c_t[1067],s_t[1067]);
fa fau_0_1068(a_i_c[1068],a_i_s[1068],b_i_c[1068],c_t[1068],s_t[1068]);
fa fau_0_1069(a_i_c[1069],a_i_s[1069],b_i_c[1069],c_t[1069],s_t[1069]);
fa fau_0_1070(a_i_c[1070],a_i_s[1070],b_i_c[1070],c_t[1070],s_t[1070]);
fa fau_0_1071(a_i_c[1071],a_i_s[1071],b_i_c[1071],c_t[1071],s_t[1071]);
fa fau_0_1072(a_i_c[1072],a_i_s[1072],b_i_c[1072],c_t[1072],s_t[1072]);
fa fau_0_1073(a_i_c[1073],a_i_s[1073],b_i_c[1073],c_t[1073],s_t[1073]);
fa fau_0_1074(a_i_c[1074],a_i_s[1074],b_i_c[1074],c_t[1074],s_t[1074]);
fa fau_0_1075(a_i_c[1075],a_i_s[1075],b_i_c[1075],c_t[1075],s_t[1075]);
fa fau_0_1076(a_i_c[1076],a_i_s[1076],b_i_c[1076],c_t[1076],s_t[1076]);
fa fau_0_1077(a_i_c[1077],a_i_s[1077],b_i_c[1077],c_t[1077],s_t[1077]);
fa fau_0_1078(a_i_c[1078],a_i_s[1078],b_i_c[1078],c_t[1078],s_t[1078]);
fa fau_0_1079(a_i_c[1079],a_i_s[1079],b_i_c[1079],c_t[1079],s_t[1079]);
fa fau_0_1080(a_i_c[1080],a_i_s[1080],b_i_c[1080],c_t[1080],s_t[1080]);
fa fau_0_1081(a_i_c[1081],a_i_s[1081],b_i_c[1081],c_t[1081],s_t[1081]);
fa fau_0_1082(a_i_c[1082],a_i_s[1082],b_i_c[1082],c_t[1082],s_t[1082]);
fa fau_0_1083(a_i_c[1083],a_i_s[1083],b_i_c[1083],c_t[1083],s_t[1083]);
fa fau_0_1084(a_i_c[1084],a_i_s[1084],b_i_c[1084],c_t[1084],s_t[1084]);
fa fau_0_1085(a_i_c[1085],a_i_s[1085],b_i_c[1085],c_t[1085],s_t[1085]);
fa fau_0_1086(a_i_c[1086],a_i_s[1086],b_i_c[1086],c_t[1086],s_t[1086]);
fa fau_0_1087(a_i_c[1087],a_i_s[1087],b_i_c[1087],c_t[1087],s_t[1087]);
fa fau_0_1088(a_i_c[1088],a_i_s[1088],b_i_c[1088],c_t[1088],s_t[1088]);
fa fau_0_1089(a_i_c[1089],a_i_s[1089],b_i_c[1089],c_t[1089],s_t[1089]);
fa fau_0_1090(a_i_c[1090],a_i_s[1090],b_i_c[1090],c_t[1090],s_t[1090]);
fa fau_0_1091(a_i_c[1091],a_i_s[1091],b_i_c[1091],c_t[1091],s_t[1091]);
fa fau_0_1092(a_i_c[1092],a_i_s[1092],b_i_c[1092],c_t[1092],s_t[1092]);
fa fau_0_1093(a_i_c[1093],a_i_s[1093],b_i_c[1093],c_t[1093],s_t[1093]);
fa fau_0_1094(a_i_c[1094],a_i_s[1094],b_i_c[1094],c_t[1094],s_t[1094]);
fa fau_0_1095(a_i_c[1095],a_i_s[1095],b_i_c[1095],c_t[1095],s_t[1095]);
fa fau_0_1096(a_i_c[1096],a_i_s[1096],b_i_c[1096],c_t[1096],s_t[1096]);
fa fau_0_1097(a_i_c[1097],a_i_s[1097],b_i_c[1097],c_t[1097],s_t[1097]);
fa fau_0_1098(a_i_c[1098],a_i_s[1098],b_i_c[1098],c_t[1098],s_t[1098]);
fa fau_0_1099(a_i_c[1099],a_i_s[1099],b_i_c[1099],c_t[1099],s_t[1099]);
fa fau_0_1100(a_i_c[1100],a_i_s[1100],b_i_c[1100],c_t[1100],s_t[1100]);
fa fau_0_1101(a_i_c[1101],a_i_s[1101],b_i_c[1101],c_t[1101],s_t[1101]);
fa fau_0_1102(a_i_c[1102],a_i_s[1102],b_i_c[1102],c_t[1102],s_t[1102]);
fa fau_0_1103(a_i_c[1103],a_i_s[1103],b_i_c[1103],c_t[1103],s_t[1103]);
fa fau_0_1104(a_i_c[1104],a_i_s[1104],b_i_c[1104],c_t[1104],s_t[1104]);
fa fau_0_1105(a_i_c[1105],a_i_s[1105],b_i_c[1105],c_t[1105],s_t[1105]);
fa fau_0_1106(a_i_c[1106],a_i_s[1106],b_i_c[1106],c_t[1106],s_t[1106]);
fa fau_0_1107(a_i_c[1107],a_i_s[1107],b_i_c[1107],c_t[1107],s_t[1107]);
fa fau_0_1108(a_i_c[1108],a_i_s[1108],b_i_c[1108],c_t[1108],s_t[1108]);
fa fau_0_1109(a_i_c[1109],a_i_s[1109],b_i_c[1109],c_t[1109],s_t[1109]);
fa fau_0_1110(a_i_c[1110],a_i_s[1110],b_i_c[1110],c_t[1110],s_t[1110]);
fa fau_0_1111(a_i_c[1111],a_i_s[1111],b_i_c[1111],c_t[1111],s_t[1111]);
fa fau_0_1112(a_i_c[1112],a_i_s[1112],b_i_c[1112],c_t[1112],s_t[1112]);
fa fau_0_1113(a_i_c[1113],a_i_s[1113],b_i_c[1113],c_t[1113],s_t[1113]);
fa fau_0_1114(a_i_c[1114],a_i_s[1114],b_i_c[1114],c_t[1114],s_t[1114]);
fa fau_0_1115(a_i_c[1115],a_i_s[1115],b_i_c[1115],c_t[1115],s_t[1115]);
fa fau_0_1116(a_i_c[1116],a_i_s[1116],b_i_c[1116],c_t[1116],s_t[1116]);
fa fau_0_1117(a_i_c[1117],a_i_s[1117],b_i_c[1117],c_t[1117],s_t[1117]);
fa fau_0_1118(a_i_c[1118],a_i_s[1118],b_i_c[1118],c_t[1118],s_t[1118]);
fa fau_0_1119(a_i_c[1119],a_i_s[1119],b_i_c[1119],c_t[1119],s_t[1119]);
fa fau_0_1120(a_i_c[1120],a_i_s[1120],b_i_c[1120],c_t[1120],s_t[1120]);
fa fau_0_1121(a_i_c[1121],a_i_s[1121],b_i_c[1121],c_t[1121],s_t[1121]);
fa fau_0_1122(a_i_c[1122],a_i_s[1122],b_i_c[1122],c_t[1122],s_t[1122]);
fa fau_0_1123(a_i_c[1123],a_i_s[1123],b_i_c[1123],c_t[1123],s_t[1123]);
fa fau_0_1124(a_i_c[1124],a_i_s[1124],b_i_c[1124],c_t[1124],s_t[1124]);
fa fau_0_1125(a_i_c[1125],a_i_s[1125],b_i_c[1125],c_t[1125],s_t[1125]);
fa fau_0_1126(a_i_c[1126],a_i_s[1126],b_i_c[1126],c_t[1126],s_t[1126]);
fa fau_0_1127(a_i_c[1127],a_i_s[1127],b_i_c[1127],c_t[1127],s_t[1127]);
fa fau_0_1128(a_i_c[1128],a_i_s[1128],b_i_c[1128],c_t[1128],s_t[1128]);
fa fau_0_1129(a_i_c[1129],a_i_s[1129],b_i_c[1129],c_t[1129],s_t[1129]);
fa fau_0_1130(a_i_c[1130],a_i_s[1130],b_i_c[1130],c_t[1130],s_t[1130]);
fa fau_0_1131(a_i_c[1131],a_i_s[1131],b_i_c[1131],c_t[1131],s_t[1131]);
fa fau_0_1132(a_i_c[1132],a_i_s[1132],b_i_c[1132],c_t[1132],s_t[1132]);
fa fau_0_1133(a_i_c[1133],a_i_s[1133],b_i_c[1133],c_t[1133],s_t[1133]);
fa fau_0_1134(a_i_c[1134],a_i_s[1134],b_i_c[1134],c_t[1134],s_t[1134]);
fa fau_0_1135(a_i_c[1135],a_i_s[1135],b_i_c[1135],c_t[1135],s_t[1135]);
fa fau_0_1136(a_i_c[1136],a_i_s[1136],b_i_c[1136],c_t[1136],s_t[1136]);
fa fau_0_1137(a_i_c[1137],a_i_s[1137],b_i_c[1137],c_t[1137],s_t[1137]);
fa fau_0_1138(a_i_c[1138],a_i_s[1138],b_i_c[1138],c_t[1138],s_t[1138]);
fa fau_0_1139(a_i_c[1139],a_i_s[1139],b_i_c[1139],c_t[1139],s_t[1139]);
fa fau_0_1140(a_i_c[1140],a_i_s[1140],b_i_c[1140],c_t[1140],s_t[1140]);
fa fau_0_1141(a_i_c[1141],a_i_s[1141],b_i_c[1141],c_t[1141],s_t[1141]);
fa fau_0_1142(a_i_c[1142],a_i_s[1142],b_i_c[1142],c_t[1142],s_t[1142]);
fa fau_0_1143(a_i_c[1143],a_i_s[1143],b_i_c[1143],c_t[1143],s_t[1143]);
fa fau_0_1144(a_i_c[1144],a_i_s[1144],b_i_c[1144],c_t[1144],s_t[1144]);
fa fau_0_1145(a_i_c[1145],a_i_s[1145],b_i_c[1145],c_t[1145],s_t[1145]);
fa fau_0_1146(a_i_c[1146],a_i_s[1146],b_i_c[1146],c_t[1146],s_t[1146]);
fa fau_0_1147(a_i_c[1147],a_i_s[1147],b_i_c[1147],c_t[1147],s_t[1147]);
fa fau_0_1148(a_i_c[1148],a_i_s[1148],b_i_c[1148],c_t[1148],s_t[1148]);
fa fau_0_1149(a_i_c[1149],a_i_s[1149],b_i_c[1149],c_t[1149],s_t[1149]);
fa fau_0_1150(a_i_c[1150],a_i_s[1150],b_i_c[1150],c_t[1150],s_t[1150]);
fa fau_0_1151(a_i_c[1151],a_i_s[1151],b_i_c[1151],c_t[1151],s_t[1151]);
fa fau_0_1152(a_i_c[1152],a_i_s[1152],b_i_c[1152],c_t[1152],s_t[1152]);
fa fau_0_1153(a_i_c[1153],a_i_s[1153],b_i_c[1153],c_t[1153],s_t[1153]);
fa fau_0_1154(a_i_c[1154],a_i_s[1154],b_i_c[1154],c_t[1154],s_t[1154]);
fa fau_0_1155(a_i_c[1155],a_i_s[1155],b_i_c[1155],c_t[1155],s_t[1155]);
fa fau_0_1156(a_i_c[1156],a_i_s[1156],b_i_c[1156],c_t[1156],s_t[1156]);
fa fau_0_1157(a_i_c[1157],a_i_s[1157],b_i_c[1157],c_t[1157],s_t[1157]);
fa fau_0_1158(a_i_c[1158],a_i_s[1158],b_i_c[1158],c_t[1158],s_t[1158]);
fa fau_0_1159(a_i_c[1159],a_i_s[1159],b_i_c[1159],c_t[1159],s_t[1159]);
fa fau_0_1160(a_i_c[1160],a_i_s[1160],b_i_c[1160],c_t[1160],s_t[1160]);
fa fau_0_1161(a_i_c[1161],a_i_s[1161],b_i_c[1161],c_t[1161],s_t[1161]);
fa fau_0_1162(a_i_c[1162],a_i_s[1162],b_i_c[1162],c_t[1162],s_t[1162]);
fa fau_0_1163(a_i_c[1163],a_i_s[1163],b_i_c[1163],c_t[1163],s_t[1163]);
fa fau_0_1164(a_i_c[1164],a_i_s[1164],b_i_c[1164],c_t[1164],s_t[1164]);
fa fau_0_1165(a_i_c[1165],a_i_s[1165],b_i_c[1165],c_t[1165],s_t[1165]);
fa fau_0_1166(a_i_c[1166],a_i_s[1166],b_i_c[1166],c_t[1166],s_t[1166]);
fa fau_0_1167(a_i_c[1167],a_i_s[1167],b_i_c[1167],c_t[1167],s_t[1167]);
fa fau_0_1168(a_i_c[1168],a_i_s[1168],b_i_c[1168],c_t[1168],s_t[1168]);
fa fau_0_1169(a_i_c[1169],a_i_s[1169],b_i_c[1169],c_t[1169],s_t[1169]);
fa fau_0_1170(a_i_c[1170],a_i_s[1170],b_i_c[1170],c_t[1170],s_t[1170]);
fa fau_0_1171(a_i_c[1171],a_i_s[1171],b_i_c[1171],c_t[1171],s_t[1171]);
fa fau_0_1172(a_i_c[1172],a_i_s[1172],b_i_c[1172],c_t[1172],s_t[1172]);
fa fau_0_1173(a_i_c[1173],a_i_s[1173],b_i_c[1173],c_t[1173],s_t[1173]);
fa fau_0_1174(a_i_c[1174],a_i_s[1174],b_i_c[1174],c_t[1174],s_t[1174]);
fa fau_0_1175(a_i_c[1175],a_i_s[1175],b_i_c[1175],c_t[1175],s_t[1175]);
fa fau_0_1176(a_i_c[1176],a_i_s[1176],b_i_c[1176],c_t[1176],s_t[1176]);
fa fau_0_1177(a_i_c[1177],a_i_s[1177],b_i_c[1177],c_t[1177],s_t[1177]);
fa fau_0_1178(a_i_c[1178],a_i_s[1178],b_i_c[1178],c_t[1178],s_t[1178]);
fa fau_0_1179(a_i_c[1179],a_i_s[1179],b_i_c[1179],c_t[1179],s_t[1179]);
fa fau_0_1180(a_i_c[1180],a_i_s[1180],b_i_c[1180],c_t[1180],s_t[1180]);
fa fau_0_1181(a_i_c[1181],a_i_s[1181],b_i_c[1181],c_t[1181],s_t[1181]);
fa fau_0_1182(a_i_c[1182],a_i_s[1182],b_i_c[1182],c_t[1182],s_t[1182]);
fa fau_0_1183(a_i_c[1183],a_i_s[1183],b_i_c[1183],c_t[1183],s_t[1183]);
fa fau_0_1184(a_i_c[1184],a_i_s[1184],b_i_c[1184],c_t[1184],s_t[1184]);
fa fau_0_1185(a_i_c[1185],a_i_s[1185],b_i_c[1185],c_t[1185],s_t[1185]);
fa fau_0_1186(a_i_c[1186],a_i_s[1186],b_i_c[1186],c_t[1186],s_t[1186]);
fa fau_0_1187(a_i_c[1187],a_i_s[1187],b_i_c[1187],c_t[1187],s_t[1187]);
fa fau_0_1188(a_i_c[1188],a_i_s[1188],b_i_c[1188],c_t[1188],s_t[1188]);
fa fau_0_1189(a_i_c[1189],a_i_s[1189],b_i_c[1189],c_t[1189],s_t[1189]);
fa fau_0_1190(a_i_c[1190],a_i_s[1190],b_i_c[1190],c_t[1190],s_t[1190]);
fa fau_0_1191(a_i_c[1191],a_i_s[1191],b_i_c[1191],c_t[1191],s_t[1191]);
fa fau_0_1192(a_i_c[1192],a_i_s[1192],b_i_c[1192],c_t[1192],s_t[1192]);
fa fau_0_1193(a_i_c[1193],a_i_s[1193],b_i_c[1193],c_t[1193],s_t[1193]);
fa fau_0_1194(a_i_c[1194],a_i_s[1194],b_i_c[1194],c_t[1194],s_t[1194]);
fa fau_0_1195(a_i_c[1195],a_i_s[1195],b_i_c[1195],c_t[1195],s_t[1195]);
fa fau_0_1196(a_i_c[1196],a_i_s[1196],b_i_c[1196],c_t[1196],s_t[1196]);
fa fau_0_1197(a_i_c[1197],a_i_s[1197],b_i_c[1197],c_t[1197],s_t[1197]);
fa fau_0_1198(a_i_c[1198],a_i_s[1198],b_i_c[1198],c_t[1198],s_t[1198]);
fa fau_0_1199(a_i_c[1199],a_i_s[1199],b_i_c[1199],c_t[1199],s_t[1199]);
fa fau_0_1200(a_i_c[1200],a_i_s[1200],b_i_c[1200],c_t[1200],s_t[1200]);
fa fau_0_1201(a_i_c[1201],a_i_s[1201],b_i_c[1201],c_t[1201],s_t[1201]);
fa fau_0_1202(a_i_c[1202],a_i_s[1202],b_i_c[1202],c_t[1202],s_t[1202]);
fa fau_0_1203(a_i_c[1203],a_i_s[1203],b_i_c[1203],c_t[1203],s_t[1203]);
fa fau_0_1204(a_i_c[1204],a_i_s[1204],b_i_c[1204],c_t[1204],s_t[1204]);
fa fau_0_1205(a_i_c[1205],a_i_s[1205],b_i_c[1205],c_t[1205],s_t[1205]);
fa fau_0_1206(a_i_c[1206],a_i_s[1206],b_i_c[1206],c_t[1206],s_t[1206]);
fa fau_0_1207(a_i_c[1207],a_i_s[1207],b_i_c[1207],c_t[1207],s_t[1207]);
fa fau_0_1208(a_i_c[1208],a_i_s[1208],b_i_c[1208],c_t[1208],s_t[1208]);
fa fau_0_1209(a_i_c[1209],a_i_s[1209],b_i_c[1209],c_t[1209],s_t[1209]);
fa fau_0_1210(a_i_c[1210],a_i_s[1210],b_i_c[1210],c_t[1210],s_t[1210]);
fa fau_0_1211(a_i_c[1211],a_i_s[1211],b_i_c[1211],c_t[1211],s_t[1211]);
fa fau_0_1212(a_i_c[1212],a_i_s[1212],b_i_c[1212],c_t[1212],s_t[1212]);
fa fau_0_1213(a_i_c[1213],a_i_s[1213],b_i_c[1213],c_t[1213],s_t[1213]);
fa fau_0_1214(a_i_c[1214],a_i_s[1214],b_i_c[1214],c_t[1214],s_t[1214]);
fa fau_0_1215(a_i_c[1215],a_i_s[1215],b_i_c[1215],c_t[1215],s_t[1215]);
fa fau_0_1216(a_i_c[1216],a_i_s[1216],b_i_c[1216],c_t[1216],s_t[1216]);
fa fau_0_1217(a_i_c[1217],a_i_s[1217],b_i_c[1217],c_t[1217],s_t[1217]);
fa fau_0_1218(a_i_c[1218],a_i_s[1218],b_i_c[1218],c_t[1218],s_t[1218]);
fa fau_0_1219(a_i_c[1219],a_i_s[1219],b_i_c[1219],c_t[1219],s_t[1219]);
fa fau_0_1220(a_i_c[1220],a_i_s[1220],b_i_c[1220],c_t[1220],s_t[1220]);
fa fau_0_1221(a_i_c[1221],a_i_s[1221],b_i_c[1221],c_t[1221],s_t[1221]);
fa fau_0_1222(a_i_c[1222],a_i_s[1222],b_i_c[1222],c_t[1222],s_t[1222]);
fa fau_0_1223(a_i_c[1223],a_i_s[1223],b_i_c[1223],c_t[1223],s_t[1223]);
fa fau_0_1224(a_i_c[1224],a_i_s[1224],b_i_c[1224],c_t[1224],s_t[1224]);
fa fau_0_1225(a_i_c[1225],a_i_s[1225],b_i_c[1225],c_t[1225],s_t[1225]);
fa fau_0_1226(a_i_c[1226],a_i_s[1226],b_i_c[1226],c_t[1226],s_t[1226]);
fa fau_0_1227(a_i_c[1227],a_i_s[1227],b_i_c[1227],c_t[1227],s_t[1227]);
fa fau_0_1228(a_i_c[1228],a_i_s[1228],b_i_c[1228],c_t[1228],s_t[1228]);
fa fau_0_1229(a_i_c[1229],a_i_s[1229],b_i_c[1229],c_t[1229],s_t[1229]);
fa fau_0_1230(a_i_c[1230],a_i_s[1230],b_i_c[1230],c_t[1230],s_t[1230]);
fa fau_0_1231(a_i_c[1231],a_i_s[1231],b_i_c[1231],c_t[1231],s_t[1231]);
fa fau_0_1232(a_i_c[1232],a_i_s[1232],b_i_c[1232],c_t[1232],s_t[1232]);
fa fau_0_1233(a_i_c[1233],a_i_s[1233],b_i_c[1233],c_t[1233],s_t[1233]);
fa fau_0_1234(a_i_c[1234],a_i_s[1234],b_i_c[1234],c_t[1234],s_t[1234]);
fa fau_0_1235(a_i_c[1235],a_i_s[1235],b_i_c[1235],c_t[1235],s_t[1235]);
fa fau_0_1236(a_i_c[1236],a_i_s[1236],b_i_c[1236],c_t[1236],s_t[1236]);
fa fau_0_1237(a_i_c[1237],a_i_s[1237],b_i_c[1237],c_t[1237],s_t[1237]);
fa fau_0_1238(a_i_c[1238],a_i_s[1238],b_i_c[1238],c_t[1238],s_t[1238]);
fa fau_0_1239(a_i_c[1239],a_i_s[1239],b_i_c[1239],c_t[1239],s_t[1239]);
fa fau_0_1240(a_i_c[1240],a_i_s[1240],b_i_c[1240],c_t[1240],s_t[1240]);
fa fau_0_1241(a_i_c[1241],a_i_s[1241],b_i_c[1241],c_t[1241],s_t[1241]);
fa fau_0_1242(a_i_c[1242],a_i_s[1242],b_i_c[1242],c_t[1242],s_t[1242]);
fa fau_0_1243(a_i_c[1243],a_i_s[1243],b_i_c[1243],c_t[1243],s_t[1243]);
fa fau_0_1244(a_i_c[1244],a_i_s[1244],b_i_c[1244],c_t[1244],s_t[1244]);
fa fau_0_1245(a_i_c[1245],a_i_s[1245],b_i_c[1245],c_t[1245],s_t[1245]);
fa fau_0_1246(a_i_c[1246],a_i_s[1246],b_i_c[1246],c_t[1246],s_t[1246]);
fa fau_0_1247(a_i_c[1247],a_i_s[1247],b_i_c[1247],c_t[1247],s_t[1247]);
fa fau_0_1248(a_i_c[1248],a_i_s[1248],b_i_c[1248],c_t[1248],s_t[1248]);
fa fau_0_1249(a_i_c[1249],a_i_s[1249],b_i_c[1249],c_t[1249],s_t[1249]);
fa fau_0_1250(a_i_c[1250],a_i_s[1250],b_i_c[1250],c_t[1250],s_t[1250]);
fa fau_0_1251(a_i_c[1251],a_i_s[1251],b_i_c[1251],c_t[1251],s_t[1251]);
fa fau_0_1252(a_i_c[1252],a_i_s[1252],b_i_c[1252],c_t[1252],s_t[1252]);
fa fau_0_1253(a_i_c[1253],a_i_s[1253],b_i_c[1253],c_t[1253],s_t[1253]);
fa fau_0_1254(a_i_c[1254],a_i_s[1254],b_i_c[1254],c_t[1254],s_t[1254]);
fa fau_0_1255(a_i_c[1255],a_i_s[1255],b_i_c[1255],c_t[1255],s_t[1255]);
fa fau_0_1256(a_i_c[1256],a_i_s[1256],b_i_c[1256],c_t[1256],s_t[1256]);
fa fau_0_1257(a_i_c[1257],a_i_s[1257],b_i_c[1257],c_t[1257],s_t[1257]);
fa fau_0_1258(a_i_c[1258],a_i_s[1258],b_i_c[1258],c_t[1258],s_t[1258]);
fa fau_0_1259(a_i_c[1259],a_i_s[1259],b_i_c[1259],c_t[1259],s_t[1259]);
fa fau_0_1260(a_i_c[1260],a_i_s[1260],b_i_c[1260],c_t[1260],s_t[1260]);
fa fau_0_1261(a_i_c[1261],a_i_s[1261],b_i_c[1261],c_t[1261],s_t[1261]);
fa fau_0_1262(a_i_c[1262],a_i_s[1262],b_i_c[1262],c_t[1262],s_t[1262]);
fa fau_0_1263(a_i_c[1263],a_i_s[1263],b_i_c[1263],c_t[1263],s_t[1263]);
fa fau_0_1264(a_i_c[1264],a_i_s[1264],b_i_c[1264],c_t[1264],s_t[1264]);
fa fau_0_1265(a_i_c[1265],a_i_s[1265],b_i_c[1265],c_t[1265],s_t[1265]);
fa fau_0_1266(a_i_c[1266],a_i_s[1266],b_i_c[1266],c_t[1266],s_t[1266]);
fa fau_0_1267(a_i_c[1267],a_i_s[1267],b_i_c[1267],c_t[1267],s_t[1267]);
fa fau_0_1268(a_i_c[1268],a_i_s[1268],b_i_c[1268],c_t[1268],s_t[1268]);
fa fau_0_1269(a_i_c[1269],a_i_s[1269],b_i_c[1269],c_t[1269],s_t[1269]);
fa fau_0_1270(a_i_c[1270],a_i_s[1270],b_i_c[1270],c_t[1270],s_t[1270]);
fa fau_0_1271(a_i_c[1271],a_i_s[1271],b_i_c[1271],c_t[1271],s_t[1271]);
fa fau_0_1272(a_i_c[1272],a_i_s[1272],b_i_c[1272],c_t[1272],s_t[1272]);
fa fau_0_1273(a_i_c[1273],a_i_s[1273],b_i_c[1273],c_t[1273],s_t[1273]);
fa fau_0_1274(a_i_c[1274],a_i_s[1274],b_i_c[1274],c_t[1274],s_t[1274]);
fa fau_0_1275(a_i_c[1275],a_i_s[1275],b_i_c[1275],c_t[1275],s_t[1275]);
fa fau_0_1276(a_i_c[1276],a_i_s[1276],b_i_c[1276],c_t[1276],s_t[1276]);
fa fau_0_1277(a_i_c[1277],a_i_s[1277],b_i_c[1277],c_t[1277],s_t[1277]);
fa fau_0_1278(a_i_c[1278],a_i_s[1278],b_i_c[1278],c_t[1278],s_t[1278]);
fa fau_0_1279(a_i_c[1279],a_i_s[1279],b_i_c[1279],c_t[1279],s_t[1279]);
fa fau_0_1280(a_i_c[1280],a_i_s[1280],b_i_c[1280],c_t[1280],s_t[1280]);
fa fau_0_1281(a_i_c[1281],a_i_s[1281],b_i_c[1281],c_t[1281],s_t[1281]);
fa fau_0_1282(a_i_c[1282],a_i_s[1282],b_i_c[1282],c_t[1282],s_t[1282]);
fa fau_0_1283(a_i_c[1283],a_i_s[1283],b_i_c[1283],c_t[1283],s_t[1283]);
fa fau_0_1284(a_i_c[1284],a_i_s[1284],b_i_c[1284],c_t[1284],s_t[1284]);
fa fau_0_1285(a_i_c[1285],a_i_s[1285],b_i_c[1285],c_t[1285],s_t[1285]);
fa fau_0_1286(a_i_c[1286],a_i_s[1286],b_i_c[1286],c_t[1286],s_t[1286]);
fa fau_0_1287(a_i_c[1287],a_i_s[1287],b_i_c[1287],c_t[1287],s_t[1287]);
fa fau_0_1288(a_i_c[1288],a_i_s[1288],b_i_c[1288],c_t[1288],s_t[1288]);
fa fau_0_1289(a_i_c[1289],a_i_s[1289],b_i_c[1289],c_t[1289],s_t[1289]);
fa fau_0_1290(a_i_c[1290],a_i_s[1290],b_i_c[1290],c_t[1290],s_t[1290]);
fa fau_0_1291(a_i_c[1291],a_i_s[1291],b_i_c[1291],c_t[1291],s_t[1291]);
fa fau_0_1292(a_i_c[1292],a_i_s[1292],b_i_c[1292],c_t[1292],s_t[1292]);
fa fau_0_1293(a_i_c[1293],a_i_s[1293],b_i_c[1293],c_t[1293],s_t[1293]);
fa fau_0_1294(a_i_c[1294],a_i_s[1294],b_i_c[1294],c_t[1294],s_t[1294]);
fa fau_0_1295(a_i_c[1295],a_i_s[1295],b_i_c[1295],c_t[1295],s_t[1295]);
fa fau_0_1296(a_i_c[1296],a_i_s[1296],b_i_c[1296],c_t[1296],s_t[1296]);
fa fau_0_1297(a_i_c[1297],a_i_s[1297],b_i_c[1297],c_t[1297],s_t[1297]);
fa fau_0_1298(a_i_c[1298],a_i_s[1298],b_i_c[1298],c_t[1298],s_t[1298]);
fa fau_0_1299(a_i_c[1299],a_i_s[1299],b_i_c[1299],c_t[1299],s_t[1299]);
fa fau_0_1300(a_i_c[1300],a_i_s[1300],b_i_c[1300],c_t[1300],s_t[1300]);
fa fau_0_1301(a_i_c[1301],a_i_s[1301],b_i_c[1301],c_t[1301],s_t[1301]);
fa fau_0_1302(a_i_c[1302],a_i_s[1302],b_i_c[1302],c_t[1302],s_t[1302]);
fa fau_0_1303(a_i_c[1303],a_i_s[1303],b_i_c[1303],c_t[1303],s_t[1303]);
fa fau_0_1304(a_i_c[1304],a_i_s[1304],b_i_c[1304],c_t[1304],s_t[1304]);
fa fau_0_1305(a_i_c[1305],a_i_s[1305],b_i_c[1305],c_t[1305],s_t[1305]);
fa fau_0_1306(a_i_c[1306],a_i_s[1306],b_i_c[1306],c_t[1306],s_t[1306]);
fa fau_0_1307(a_i_c[1307],a_i_s[1307],b_i_c[1307],c_t[1307],s_t[1307]);
fa fau_0_1308(a_i_c[1308],a_i_s[1308],b_i_c[1308],c_t[1308],s_t[1308]);
fa fau_0_1309(a_i_c[1309],a_i_s[1309],b_i_c[1309],c_t[1309],s_t[1309]);
fa fau_0_1310(a_i_c[1310],a_i_s[1310],b_i_c[1310],c_t[1310],s_t[1310]);
fa fau_0_1311(a_i_c[1311],a_i_s[1311],b_i_c[1311],c_t[1311],s_t[1311]);
fa fau_0_1312(a_i_c[1312],a_i_s[1312],b_i_c[1312],c_t[1312],s_t[1312]);
fa fau_0_1313(a_i_c[1313],a_i_s[1313],b_i_c[1313],c_t[1313],s_t[1313]);
fa fau_0_1314(a_i_c[1314],a_i_s[1314],b_i_c[1314],c_t[1314],s_t[1314]);
fa fau_0_1315(a_i_c[1315],a_i_s[1315],b_i_c[1315],c_t[1315],s_t[1315]);
fa fau_0_1316(a_i_c[1316],a_i_s[1316],b_i_c[1316],c_t[1316],s_t[1316]);
fa fau_0_1317(a_i_c[1317],a_i_s[1317],b_i_c[1317],c_t[1317],s_t[1317]);
fa fau_0_1318(a_i_c[1318],a_i_s[1318],b_i_c[1318],c_t[1318],s_t[1318]);
fa fau_0_1319(a_i_c[1319],a_i_s[1319],b_i_c[1319],c_t[1319],s_t[1319]);
fa fau_0_1320(a_i_c[1320],a_i_s[1320],b_i_c[1320],c_t[1320],s_t[1320]);
fa fau_0_1321(a_i_c[1321],a_i_s[1321],b_i_c[1321],c_t[1321],s_t[1321]);
fa fau_0_1322(a_i_c[1322],a_i_s[1322],b_i_c[1322],c_t[1322],s_t[1322]);
fa fau_0_1323(a_i_c[1323],a_i_s[1323],b_i_c[1323],c_t[1323],s_t[1323]);
fa fau_0_1324(a_i_c[1324],a_i_s[1324],b_i_c[1324],c_t[1324],s_t[1324]);
fa fau_0_1325(a_i_c[1325],a_i_s[1325],b_i_c[1325],c_t[1325],s_t[1325]);
fa fau_0_1326(a_i_c[1326],a_i_s[1326],b_i_c[1326],c_t[1326],s_t[1326]);
fa fau_0_1327(a_i_c[1327],a_i_s[1327],b_i_c[1327],c_t[1327],s_t[1327]);
fa fau_0_1328(a_i_c[1328],a_i_s[1328],b_i_c[1328],c_t[1328],s_t[1328]);
fa fau_0_1329(a_i_c[1329],a_i_s[1329],b_i_c[1329],c_t[1329],s_t[1329]);
fa fau_0_1330(a_i_c[1330],a_i_s[1330],b_i_c[1330],c_t[1330],s_t[1330]);
fa fau_0_1331(a_i_c[1331],a_i_s[1331],b_i_c[1331],c_t[1331],s_t[1331]);
fa fau_0_1332(a_i_c[1332],a_i_s[1332],b_i_c[1332],c_t[1332],s_t[1332]);
fa fau_0_1333(a_i_c[1333],a_i_s[1333],b_i_c[1333],c_t[1333],s_t[1333]);
fa fau_0_1334(a_i_c[1334],a_i_s[1334],b_i_c[1334],c_t[1334],s_t[1334]);
fa fau_0_1335(a_i_c[1335],a_i_s[1335],b_i_c[1335],c_t[1335],s_t[1335]);
fa fau_0_1336(a_i_c[1336],a_i_s[1336],b_i_c[1336],c_t[1336],s_t[1336]);
fa fau_0_1337(a_i_c[1337],a_i_s[1337],b_i_c[1337],c_t[1337],s_t[1337]);
fa fau_0_1338(a_i_c[1338],a_i_s[1338],b_i_c[1338],c_t[1338],s_t[1338]);
fa fau_0_1339(a_i_c[1339],a_i_s[1339],b_i_c[1339],c_t[1339],s_t[1339]);
fa fau_0_1340(a_i_c[1340],a_i_s[1340],b_i_c[1340],c_t[1340],s_t[1340]);
fa fau_0_1341(a_i_c[1341],a_i_s[1341],b_i_c[1341],c_t[1341],s_t[1341]);
fa fau_0_1342(a_i_c[1342],a_i_s[1342],b_i_c[1342],c_t[1342],s_t[1342]);
fa fau_0_1343(a_i_c[1343],a_i_s[1343],b_i_c[1343],c_t[1343],s_t[1343]);
fa fau_0_1344(a_i_c[1344],a_i_s[1344],b_i_c[1344],c_t[1344],s_t[1344]);
fa fau_0_1345(a_i_c[1345],a_i_s[1345],b_i_c[1345],c_t[1345],s_t[1345]);
fa fau_0_1346(a_i_c[1346],a_i_s[1346],b_i_c[1346],c_t[1346],s_t[1346]);
fa fau_0_1347(a_i_c[1347],a_i_s[1347],b_i_c[1347],c_t[1347],s_t[1347]);
fa fau_0_1348(a_i_c[1348],a_i_s[1348],b_i_c[1348],c_t[1348],s_t[1348]);
fa fau_0_1349(a_i_c[1349],a_i_s[1349],b_i_c[1349],c_t[1349],s_t[1349]);
fa fau_0_1350(a_i_c[1350],a_i_s[1350],b_i_c[1350],c_t[1350],s_t[1350]);
fa fau_0_1351(a_i_c[1351],a_i_s[1351],b_i_c[1351],c_t[1351],s_t[1351]);
fa fau_0_1352(a_i_c[1352],a_i_s[1352],b_i_c[1352],c_t[1352],s_t[1352]);
fa fau_0_1353(a_i_c[1353],a_i_s[1353],b_i_c[1353],c_t[1353],s_t[1353]);
fa fau_0_1354(a_i_c[1354],a_i_s[1354],b_i_c[1354],c_t[1354],s_t[1354]);
fa fau_0_1355(a_i_c[1355],a_i_s[1355],b_i_c[1355],c_t[1355],s_t[1355]);
fa fau_0_1356(a_i_c[1356],a_i_s[1356],b_i_c[1356],c_t[1356],s_t[1356]);
fa fau_0_1357(a_i_c[1357],a_i_s[1357],b_i_c[1357],c_t[1357],s_t[1357]);
fa fau_0_1358(a_i_c[1358],a_i_s[1358],b_i_c[1358],c_t[1358],s_t[1358]);
fa fau_0_1359(a_i_c[1359],a_i_s[1359],b_i_c[1359],c_t[1359],s_t[1359]);
fa fau_0_1360(a_i_c[1360],a_i_s[1360],b_i_c[1360],c_t[1360],s_t[1360]);
fa fau_0_1361(a_i_c[1361],a_i_s[1361],b_i_c[1361],c_t[1361],s_t[1361]);
fa fau_0_1362(a_i_c[1362],a_i_s[1362],b_i_c[1362],c_t[1362],s_t[1362]);
fa fau_0_1363(a_i_c[1363],a_i_s[1363],b_i_c[1363],c_t[1363],s_t[1363]);
fa fau_0_1364(a_i_c[1364],a_i_s[1364],b_i_c[1364],c_t[1364],s_t[1364]);
fa fau_0_1365(a_i_c[1365],a_i_s[1365],b_i_c[1365],c_t[1365],s_t[1365]);
fa fau_0_1366(a_i_c[1366],a_i_s[1366],b_i_c[1366],c_t[1366],s_t[1366]);
fa fau_0_1367(a_i_c[1367],a_i_s[1367],b_i_c[1367],c_t[1367],s_t[1367]);
fa fau_0_1368(a_i_c[1368],a_i_s[1368],b_i_c[1368],c_t[1368],s_t[1368]);
fa fau_0_1369(a_i_c[1369],a_i_s[1369],b_i_c[1369],c_t[1369],s_t[1369]);
fa fau_0_1370(a_i_c[1370],a_i_s[1370],b_i_c[1370],c_t[1370],s_t[1370]);
fa fau_0_1371(a_i_c[1371],a_i_s[1371],b_i_c[1371],c_t[1371],s_t[1371]);
fa fau_0_1372(a_i_c[1372],a_i_s[1372],b_i_c[1372],c_t[1372],s_t[1372]);
fa fau_0_1373(a_i_c[1373],a_i_s[1373],b_i_c[1373],c_t[1373],s_t[1373]);
fa fau_0_1374(a_i_c[1374],a_i_s[1374],b_i_c[1374],c_t[1374],s_t[1374]);
fa fau_0_1375(a_i_c[1375],a_i_s[1375],b_i_c[1375],c_t[1375],s_t[1375]);
fa fau_0_1376(a_i_c[1376],a_i_s[1376],b_i_c[1376],c_t[1376],s_t[1376]);
fa fau_0_1377(a_i_c[1377],a_i_s[1377],b_i_c[1377],c_t[1377],s_t[1377]);
fa fau_0_1378(a_i_c[1378],a_i_s[1378],b_i_c[1378],c_t[1378],s_t[1378]);
fa fau_0_1379(a_i_c[1379],a_i_s[1379],b_i_c[1379],c_t[1379],s_t[1379]);
fa fau_0_1380(a_i_c[1380],a_i_s[1380],b_i_c[1380],c_t[1380],s_t[1380]);
fa fau_0_1381(a_i_c[1381],a_i_s[1381],b_i_c[1381],c_t[1381],s_t[1381]);
fa fau_0_1382(a_i_c[1382],a_i_s[1382],b_i_c[1382],c_t[1382],s_t[1382]);
fa fau_0_1383(a_i_c[1383],a_i_s[1383],b_i_c[1383],c_t[1383],s_t[1383]);
fa fau_0_1384(a_i_c[1384],a_i_s[1384],b_i_c[1384],c_t[1384],s_t[1384]);
fa fau_0_1385(a_i_c[1385],a_i_s[1385],b_i_c[1385],c_t[1385],s_t[1385]);
fa fau_0_1386(a_i_c[1386],a_i_s[1386],b_i_c[1386],c_t[1386],s_t[1386]);
fa fau_0_1387(a_i_c[1387],a_i_s[1387],b_i_c[1387],c_t[1387],s_t[1387]);
fa fau_0_1388(a_i_c[1388],a_i_s[1388],b_i_c[1388],c_t[1388],s_t[1388]);
fa fau_0_1389(a_i_c[1389],a_i_s[1389],b_i_c[1389],c_t[1389],s_t[1389]);
fa fau_0_1390(a_i_c[1390],a_i_s[1390],b_i_c[1390],c_t[1390],s_t[1390]);
fa fau_0_1391(a_i_c[1391],a_i_s[1391],b_i_c[1391],c_t[1391],s_t[1391]);
fa fau_0_1392(a_i_c[1392],a_i_s[1392],b_i_c[1392],c_t[1392],s_t[1392]);
fa fau_0_1393(a_i_c[1393],a_i_s[1393],b_i_c[1393],c_t[1393],s_t[1393]);
fa fau_0_1394(a_i_c[1394],a_i_s[1394],b_i_c[1394],c_t[1394],s_t[1394]);
fa fau_0_1395(a_i_c[1395],a_i_s[1395],b_i_c[1395],c_t[1395],s_t[1395]);
fa fau_0_1396(a_i_c[1396],a_i_s[1396],b_i_c[1396],c_t[1396],s_t[1396]);
fa fau_0_1397(a_i_c[1397],a_i_s[1397],b_i_c[1397],c_t[1397],s_t[1397]);
fa fau_0_1398(a_i_c[1398],a_i_s[1398],b_i_c[1398],c_t[1398],s_t[1398]);
fa fau_0_1399(a_i_c[1399],a_i_s[1399],b_i_c[1399],c_t[1399],s_t[1399]);
fa fau_0_1400(a_i_c[1400],a_i_s[1400],b_i_c[1400],c_t[1400],s_t[1400]);
fa fau_0_1401(a_i_c[1401],a_i_s[1401],b_i_c[1401],c_t[1401],s_t[1401]);
fa fau_0_1402(a_i_c[1402],a_i_s[1402],b_i_c[1402],c_t[1402],s_t[1402]);
fa fau_0_1403(a_i_c[1403],a_i_s[1403],b_i_c[1403],c_t[1403],s_t[1403]);
fa fau_0_1404(a_i_c[1404],a_i_s[1404],b_i_c[1404],c_t[1404],s_t[1404]);
fa fau_0_1405(a_i_c[1405],a_i_s[1405],b_i_c[1405],c_t[1405],s_t[1405]);
fa fau_0_1406(a_i_c[1406],a_i_s[1406],b_i_c[1406],c_t[1406],s_t[1406]);
fa fau_0_1407(a_i_c[1407],a_i_s[1407],b_i_c[1407],c_t[1407],s_t[1407]);
fa fau_0_1408(a_i_c[1408],a_i_s[1408],b_i_c[1408],c_t[1408],s_t[1408]);
fa fau_0_1409(a_i_c[1409],a_i_s[1409],b_i_c[1409],c_t[1409],s_t[1409]);
fa fau_0_1410(a_i_c[1410],a_i_s[1410],b_i_c[1410],c_t[1410],s_t[1410]);
fa fau_0_1411(a_i_c[1411],a_i_s[1411],b_i_c[1411],c_t[1411],s_t[1411]);
fa fau_0_1412(a_i_c[1412],a_i_s[1412],b_i_c[1412],c_t[1412],s_t[1412]);
fa fau_0_1413(a_i_c[1413],a_i_s[1413],b_i_c[1413],c_t[1413],s_t[1413]);
fa fau_0_1414(a_i_c[1414],a_i_s[1414],b_i_c[1414],c_t[1414],s_t[1414]);
fa fau_0_1415(a_i_c[1415],a_i_s[1415],b_i_c[1415],c_t[1415],s_t[1415]);
fa fau_0_1416(a_i_c[1416],a_i_s[1416],b_i_c[1416],c_t[1416],s_t[1416]);
fa fau_0_1417(a_i_c[1417],a_i_s[1417],b_i_c[1417],c_t[1417],s_t[1417]);
fa fau_0_1418(a_i_c[1418],a_i_s[1418],b_i_c[1418],c_t[1418],s_t[1418]);
fa fau_0_1419(a_i_c[1419],a_i_s[1419],b_i_c[1419],c_t[1419],s_t[1419]);
fa fau_0_1420(a_i_c[1420],a_i_s[1420],b_i_c[1420],c_t[1420],s_t[1420]);
fa fau_0_1421(a_i_c[1421],a_i_s[1421],b_i_c[1421],c_t[1421],s_t[1421]);
fa fau_0_1422(a_i_c[1422],a_i_s[1422],b_i_c[1422],c_t[1422],s_t[1422]);
fa fau_0_1423(a_i_c[1423],a_i_s[1423],b_i_c[1423],c_t[1423],s_t[1423]);
fa fau_0_1424(a_i_c[1424],a_i_s[1424],b_i_c[1424],c_t[1424],s_t[1424]);
fa fau_0_1425(a_i_c[1425],a_i_s[1425],b_i_c[1425],c_t[1425],s_t[1425]);
fa fau_0_1426(a_i_c[1426],a_i_s[1426],b_i_c[1426],c_t[1426],s_t[1426]);
fa fau_0_1427(a_i_c[1427],a_i_s[1427],b_i_c[1427],c_t[1427],s_t[1427]);
fa fau_0_1428(a_i_c[1428],a_i_s[1428],b_i_c[1428],c_t[1428],s_t[1428]);
fa fau_0_1429(a_i_c[1429],a_i_s[1429],b_i_c[1429],c_t[1429],s_t[1429]);
fa fau_0_1430(a_i_c[1430],a_i_s[1430],b_i_c[1430],c_t[1430],s_t[1430]);
fa fau_0_1431(a_i_c[1431],a_i_s[1431],b_i_c[1431],c_t[1431],s_t[1431]);
fa fau_0_1432(a_i_c[1432],a_i_s[1432],b_i_c[1432],c_t[1432],s_t[1432]);
fa fau_0_1433(a_i_c[1433],a_i_s[1433],b_i_c[1433],c_t[1433],s_t[1433]);
fa fau_0_1434(a_i_c[1434],a_i_s[1434],b_i_c[1434],c_t[1434],s_t[1434]);
fa fau_0_1435(a_i_c[1435],a_i_s[1435],b_i_c[1435],c_t[1435],s_t[1435]);
fa fau_0_1436(a_i_c[1436],a_i_s[1436],b_i_c[1436],c_t[1436],s_t[1436]);
fa fau_0_1437(a_i_c[1437],a_i_s[1437],b_i_c[1437],c_t[1437],s_t[1437]);
fa fau_0_1438(a_i_c[1438],a_i_s[1438],b_i_c[1438],c_t[1438],s_t[1438]);
fa fau_0_1439(a_i_c[1439],a_i_s[1439],b_i_c[1439],c_t[1439],s_t[1439]);
fa fau_0_1440(a_i_c[1440],a_i_s[1440],b_i_c[1440],c_t[1440],s_t[1440]);
fa fau_0_1441(a_i_c[1441],a_i_s[1441],b_i_c[1441],c_t[1441],s_t[1441]);
fa fau_0_1442(a_i_c[1442],a_i_s[1442],b_i_c[1442],c_t[1442],s_t[1442]);
fa fau_0_1443(a_i_c[1443],a_i_s[1443],b_i_c[1443],c_t[1443],s_t[1443]);
fa fau_0_1444(a_i_c[1444],a_i_s[1444],b_i_c[1444],c_t[1444],s_t[1444]);
fa fau_0_1445(a_i_c[1445],a_i_s[1445],b_i_c[1445],c_t[1445],s_t[1445]);
fa fau_0_1446(a_i_c[1446],a_i_s[1446],b_i_c[1446],c_t[1446],s_t[1446]);
fa fau_0_1447(a_i_c[1447],a_i_s[1447],b_i_c[1447],c_t[1447],s_t[1447]);
fa fau_0_1448(a_i_c[1448],a_i_s[1448],b_i_c[1448],c_t[1448],s_t[1448]);
fa fau_0_1449(a_i_c[1449],a_i_s[1449],b_i_c[1449],c_t[1449],s_t[1449]);
fa fau_0_1450(a_i_c[1450],a_i_s[1450],b_i_c[1450],c_t[1450],s_t[1450]);
fa fau_0_1451(a_i_c[1451],a_i_s[1451],b_i_c[1451],c_t[1451],s_t[1451]);
fa fau_0_1452(a_i_c[1452],a_i_s[1452],b_i_c[1452],c_t[1452],s_t[1452]);
fa fau_0_1453(a_i_c[1453],a_i_s[1453],b_i_c[1453],c_t[1453],s_t[1453]);
fa fau_0_1454(a_i_c[1454],a_i_s[1454],b_i_c[1454],c_t[1454],s_t[1454]);
fa fau_0_1455(a_i_c[1455],a_i_s[1455],b_i_c[1455],c_t[1455],s_t[1455]);
fa fau_0_1456(a_i_c[1456],a_i_s[1456],b_i_c[1456],c_t[1456],s_t[1456]);
fa fau_0_1457(a_i_c[1457],a_i_s[1457],b_i_c[1457],c_t[1457],s_t[1457]);
fa fau_0_1458(a_i_c[1458],a_i_s[1458],b_i_c[1458],c_t[1458],s_t[1458]);
fa fau_0_1459(a_i_c[1459],a_i_s[1459],b_i_c[1459],c_t[1459],s_t[1459]);
fa fau_0_1460(a_i_c[1460],a_i_s[1460],b_i_c[1460],c_t[1460],s_t[1460]);
fa fau_0_1461(a_i_c[1461],a_i_s[1461],b_i_c[1461],c_t[1461],s_t[1461]);
fa fau_0_1462(a_i_c[1462],a_i_s[1462],b_i_c[1462],c_t[1462],s_t[1462]);
fa fau_0_1463(a_i_c[1463],a_i_s[1463],b_i_c[1463],c_t[1463],s_t[1463]);
fa fau_0_1464(a_i_c[1464],a_i_s[1464],b_i_c[1464],c_t[1464],s_t[1464]);
fa fau_0_1465(a_i_c[1465],a_i_s[1465],b_i_c[1465],c_t[1465],s_t[1465]);
fa fau_0_1466(a_i_c[1466],a_i_s[1466],b_i_c[1466],c_t[1466],s_t[1466]);
fa fau_0_1467(a_i_c[1467],a_i_s[1467],b_i_c[1467],c_t[1467],s_t[1467]);
fa fau_0_1468(a_i_c[1468],a_i_s[1468],b_i_c[1468],c_t[1468],s_t[1468]);
fa fau_0_1469(a_i_c[1469],a_i_s[1469],b_i_c[1469],c_t[1469],s_t[1469]);
fa fau_0_1470(a_i_c[1470],a_i_s[1470],b_i_c[1470],c_t[1470],s_t[1470]);
fa fau_0_1471(a_i_c[1471],a_i_s[1471],b_i_c[1471],c_t[1471],s_t[1471]);
fa fau_0_1472(a_i_c[1472],a_i_s[1472],b_i_c[1472],c_t[1472],s_t[1472]);
fa fau_0_1473(a_i_c[1473],a_i_s[1473],b_i_c[1473],c_t[1473],s_t[1473]);
fa fau_0_1474(a_i_c[1474],a_i_s[1474],b_i_c[1474],c_t[1474],s_t[1474]);
fa fau_0_1475(a_i_c[1475],a_i_s[1475],b_i_c[1475],c_t[1475],s_t[1475]);
fa fau_0_1476(a_i_c[1476],a_i_s[1476],b_i_c[1476],c_t[1476],s_t[1476]);
fa fau_0_1477(a_i_c[1477],a_i_s[1477],b_i_c[1477],c_t[1477],s_t[1477]);
fa fau_0_1478(a_i_c[1478],a_i_s[1478],b_i_c[1478],c_t[1478],s_t[1478]);
fa fau_0_1479(a_i_c[1479],a_i_s[1479],b_i_c[1479],c_t[1479],s_t[1479]);
fa fau_0_1480(a_i_c[1480],a_i_s[1480],b_i_c[1480],c_t[1480],s_t[1480]);
fa fau_0_1481(a_i_c[1481],a_i_s[1481],b_i_c[1481],c_t[1481],s_t[1481]);
fa fau_0_1482(a_i_c[1482],a_i_s[1482],b_i_c[1482],c_t[1482],s_t[1482]);
fa fau_0_1483(a_i_c[1483],a_i_s[1483],b_i_c[1483],c_t[1483],s_t[1483]);
fa fau_0_1484(a_i_c[1484],a_i_s[1484],b_i_c[1484],c_t[1484],s_t[1484]);
fa fau_0_1485(a_i_c[1485],a_i_s[1485],b_i_c[1485],c_t[1485],s_t[1485]);
fa fau_0_1486(a_i_c[1486],a_i_s[1486],b_i_c[1486],c_t[1486],s_t[1486]);
fa fau_0_1487(a_i_c[1487],a_i_s[1487],b_i_c[1487],c_t[1487],s_t[1487]);
fa fau_0_1488(a_i_c[1488],a_i_s[1488],b_i_c[1488],c_t[1488],s_t[1488]);
fa fau_0_1489(a_i_c[1489],a_i_s[1489],b_i_c[1489],c_t[1489],s_t[1489]);
fa fau_0_1490(a_i_c[1490],a_i_s[1490],b_i_c[1490],c_t[1490],s_t[1490]);
fa fau_0_1491(a_i_c[1491],a_i_s[1491],b_i_c[1491],c_t[1491],s_t[1491]);
fa fau_0_1492(a_i_c[1492],a_i_s[1492],b_i_c[1492],c_t[1492],s_t[1492]);
fa fau_0_1493(a_i_c[1493],a_i_s[1493],b_i_c[1493],c_t[1493],s_t[1493]);
fa fau_0_1494(a_i_c[1494],a_i_s[1494],b_i_c[1494],c_t[1494],s_t[1494]);
fa fau_0_1495(a_i_c[1495],a_i_s[1495],b_i_c[1495],c_t[1495],s_t[1495]);
fa fau_0_1496(a_i_c[1496],a_i_s[1496],b_i_c[1496],c_t[1496],s_t[1496]);
fa fau_0_1497(a_i_c[1497],a_i_s[1497],b_i_c[1497],c_t[1497],s_t[1497]);
fa fau_0_1498(a_i_c[1498],a_i_s[1498],b_i_c[1498],c_t[1498],s_t[1498]);
fa fau_0_1499(a_i_c[1499],a_i_s[1499],b_i_c[1499],c_t[1499],s_t[1499]);
fa fau_0_1500(a_i_c[1500],a_i_s[1500],b_i_c[1500],c_t[1500],s_t[1500]);
fa fau_0_1501(a_i_c[1501],a_i_s[1501],b_i_c[1501],c_t[1501],s_t[1501]);
fa fau_0_1502(a_i_c[1502],a_i_s[1502],b_i_c[1502],c_t[1502],s_t[1502]);
fa fau_0_1503(a_i_c[1503],a_i_s[1503],b_i_c[1503],c_t[1503],s_t[1503]);
fa fau_0_1504(a_i_c[1504],a_i_s[1504],b_i_c[1504],c_t[1504],s_t[1504]);
fa fau_0_1505(a_i_c[1505],a_i_s[1505],b_i_c[1505],c_t[1505],s_t[1505]);
    
fa fau_1_1(b_i_s[1],s_t[1],c_t[0],c_t2[1],s_t2[1]);
fa fau_1_2(b_i_s[2],s_t[2],c_t[1],c_t2[2],s_t2[2]);
fa fau_1_3(b_i_s[3],s_t[3],c_t[2],c_t2[3],s_t2[3]);
fa fau_1_4(b_i_s[4],s_t[4],c_t[3],c_t2[4],s_t2[4]);
fa fau_1_5(b_i_s[5],s_t[5],c_t[4],c_t2[5],s_t2[5]);
fa fau_1_6(b_i_s[6],s_t[6],c_t[5],c_t2[6],s_t2[6]);
fa fau_1_7(b_i_s[7],s_t[7],c_t[6],c_t2[7],s_t2[7]);
fa fau_1_8(b_i_s[8],s_t[8],c_t[7],c_t2[8],s_t2[8]);
fa fau_1_9(b_i_s[9],s_t[9],c_t[8],c_t2[9],s_t2[9]);
fa fau_1_10(b_i_s[10],s_t[10],c_t[9],c_t2[10],s_t2[10]);
fa fau_1_11(b_i_s[11],s_t[11],c_t[10],c_t2[11],s_t2[11]);
fa fau_1_12(b_i_s[12],s_t[12],c_t[11],c_t2[12],s_t2[12]);
fa fau_1_13(b_i_s[13],s_t[13],c_t[12],c_t2[13],s_t2[13]);
fa fau_1_14(b_i_s[14],s_t[14],c_t[13],c_t2[14],s_t2[14]);
fa fau_1_15(b_i_s[15],s_t[15],c_t[14],c_t2[15],s_t2[15]);
fa fau_1_16(b_i_s[16],s_t[16],c_t[15],c_t2[16],s_t2[16]);
fa fau_1_17(b_i_s[17],s_t[17],c_t[16],c_t2[17],s_t2[17]);
fa fau_1_18(b_i_s[18],s_t[18],c_t[17],c_t2[18],s_t2[18]);
fa fau_1_19(b_i_s[19],s_t[19],c_t[18],c_t2[19],s_t2[19]);
fa fau_1_20(b_i_s[20],s_t[20],c_t[19],c_t2[20],s_t2[20]);
fa fau_1_21(b_i_s[21],s_t[21],c_t[20],c_t2[21],s_t2[21]);
fa fau_1_22(b_i_s[22],s_t[22],c_t[21],c_t2[22],s_t2[22]);
fa fau_1_23(b_i_s[23],s_t[23],c_t[22],c_t2[23],s_t2[23]);
fa fau_1_24(b_i_s[24],s_t[24],c_t[23],c_t2[24],s_t2[24]);
fa fau_1_25(b_i_s[25],s_t[25],c_t[24],c_t2[25],s_t2[25]);
fa fau_1_26(b_i_s[26],s_t[26],c_t[25],c_t2[26],s_t2[26]);
fa fau_1_27(b_i_s[27],s_t[27],c_t[26],c_t2[27],s_t2[27]);
fa fau_1_28(b_i_s[28],s_t[28],c_t[27],c_t2[28],s_t2[28]);
fa fau_1_29(b_i_s[29],s_t[29],c_t[28],c_t2[29],s_t2[29]);
fa fau_1_30(b_i_s[30],s_t[30],c_t[29],c_t2[30],s_t2[30]);
fa fau_1_31(b_i_s[31],s_t[31],c_t[30],c_t2[31],s_t2[31]);
fa fau_1_32(b_i_s[32],s_t[32],c_t[31],c_t2[32],s_t2[32]);
fa fau_1_33(b_i_s[33],s_t[33],c_t[32],c_t2[33],s_t2[33]);
fa fau_1_34(b_i_s[34],s_t[34],c_t[33],c_t2[34],s_t2[34]);
fa fau_1_35(b_i_s[35],s_t[35],c_t[34],c_t2[35],s_t2[35]);
fa fau_1_36(b_i_s[36],s_t[36],c_t[35],c_t2[36],s_t2[36]);
fa fau_1_37(b_i_s[37],s_t[37],c_t[36],c_t2[37],s_t2[37]);
fa fau_1_38(b_i_s[38],s_t[38],c_t[37],c_t2[38],s_t2[38]);
fa fau_1_39(b_i_s[39],s_t[39],c_t[38],c_t2[39],s_t2[39]);
fa fau_1_40(b_i_s[40],s_t[40],c_t[39],c_t2[40],s_t2[40]);
fa fau_1_41(b_i_s[41],s_t[41],c_t[40],c_t2[41],s_t2[41]);
fa fau_1_42(b_i_s[42],s_t[42],c_t[41],c_t2[42],s_t2[42]);
fa fau_1_43(b_i_s[43],s_t[43],c_t[42],c_t2[43],s_t2[43]);
fa fau_1_44(b_i_s[44],s_t[44],c_t[43],c_t2[44],s_t2[44]);
fa fau_1_45(b_i_s[45],s_t[45],c_t[44],c_t2[45],s_t2[45]);
fa fau_1_46(b_i_s[46],s_t[46],c_t[45],c_t2[46],s_t2[46]);
fa fau_1_47(b_i_s[47],s_t[47],c_t[46],c_t2[47],s_t2[47]);
fa fau_1_48(b_i_s[48],s_t[48],c_t[47],c_t2[48],s_t2[48]);
fa fau_1_49(b_i_s[49],s_t[49],c_t[48],c_t2[49],s_t2[49]);
fa fau_1_50(b_i_s[50],s_t[50],c_t[49],c_t2[50],s_t2[50]);
fa fau_1_51(b_i_s[51],s_t[51],c_t[50],c_t2[51],s_t2[51]);
fa fau_1_52(b_i_s[52],s_t[52],c_t[51],c_t2[52],s_t2[52]);
fa fau_1_53(b_i_s[53],s_t[53],c_t[52],c_t2[53],s_t2[53]);
fa fau_1_54(b_i_s[54],s_t[54],c_t[53],c_t2[54],s_t2[54]);
fa fau_1_55(b_i_s[55],s_t[55],c_t[54],c_t2[55],s_t2[55]);
fa fau_1_56(b_i_s[56],s_t[56],c_t[55],c_t2[56],s_t2[56]);
fa fau_1_57(b_i_s[57],s_t[57],c_t[56],c_t2[57],s_t2[57]);
fa fau_1_58(b_i_s[58],s_t[58],c_t[57],c_t2[58],s_t2[58]);
fa fau_1_59(b_i_s[59],s_t[59],c_t[58],c_t2[59],s_t2[59]);
fa fau_1_60(b_i_s[60],s_t[60],c_t[59],c_t2[60],s_t2[60]);
fa fau_1_61(b_i_s[61],s_t[61],c_t[60],c_t2[61],s_t2[61]);
fa fau_1_62(b_i_s[62],s_t[62],c_t[61],c_t2[62],s_t2[62]);
fa fau_1_63(b_i_s[63],s_t[63],c_t[62],c_t2[63],s_t2[63]);
fa fau_1_64(b_i_s[64],s_t[64],c_t[63],c_t2[64],s_t2[64]);
fa fau_1_65(b_i_s[65],s_t[65],c_t[64],c_t2[65],s_t2[65]);
fa fau_1_66(b_i_s[66],s_t[66],c_t[65],c_t2[66],s_t2[66]);
fa fau_1_67(b_i_s[67],s_t[67],c_t[66],c_t2[67],s_t2[67]);
fa fau_1_68(b_i_s[68],s_t[68],c_t[67],c_t2[68],s_t2[68]);
fa fau_1_69(b_i_s[69],s_t[69],c_t[68],c_t2[69],s_t2[69]);
fa fau_1_70(b_i_s[70],s_t[70],c_t[69],c_t2[70],s_t2[70]);
fa fau_1_71(b_i_s[71],s_t[71],c_t[70],c_t2[71],s_t2[71]);
fa fau_1_72(b_i_s[72],s_t[72],c_t[71],c_t2[72],s_t2[72]);
fa fau_1_73(b_i_s[73],s_t[73],c_t[72],c_t2[73],s_t2[73]);
fa fau_1_74(b_i_s[74],s_t[74],c_t[73],c_t2[74],s_t2[74]);
fa fau_1_75(b_i_s[75],s_t[75],c_t[74],c_t2[75],s_t2[75]);
fa fau_1_76(b_i_s[76],s_t[76],c_t[75],c_t2[76],s_t2[76]);
fa fau_1_77(b_i_s[77],s_t[77],c_t[76],c_t2[77],s_t2[77]);
fa fau_1_78(b_i_s[78],s_t[78],c_t[77],c_t2[78],s_t2[78]);
fa fau_1_79(b_i_s[79],s_t[79],c_t[78],c_t2[79],s_t2[79]);
fa fau_1_80(b_i_s[80],s_t[80],c_t[79],c_t2[80],s_t2[80]);
fa fau_1_81(b_i_s[81],s_t[81],c_t[80],c_t2[81],s_t2[81]);
fa fau_1_82(b_i_s[82],s_t[82],c_t[81],c_t2[82],s_t2[82]);
fa fau_1_83(b_i_s[83],s_t[83],c_t[82],c_t2[83],s_t2[83]);
fa fau_1_84(b_i_s[84],s_t[84],c_t[83],c_t2[84],s_t2[84]);
fa fau_1_85(b_i_s[85],s_t[85],c_t[84],c_t2[85],s_t2[85]);
fa fau_1_86(b_i_s[86],s_t[86],c_t[85],c_t2[86],s_t2[86]);
fa fau_1_87(b_i_s[87],s_t[87],c_t[86],c_t2[87],s_t2[87]);
fa fau_1_88(b_i_s[88],s_t[88],c_t[87],c_t2[88],s_t2[88]);
fa fau_1_89(b_i_s[89],s_t[89],c_t[88],c_t2[89],s_t2[89]);
fa fau_1_90(b_i_s[90],s_t[90],c_t[89],c_t2[90],s_t2[90]);
fa fau_1_91(b_i_s[91],s_t[91],c_t[90],c_t2[91],s_t2[91]);
fa fau_1_92(b_i_s[92],s_t[92],c_t[91],c_t2[92],s_t2[92]);
fa fau_1_93(b_i_s[93],s_t[93],c_t[92],c_t2[93],s_t2[93]);
fa fau_1_94(b_i_s[94],s_t[94],c_t[93],c_t2[94],s_t2[94]);
fa fau_1_95(b_i_s[95],s_t[95],c_t[94],c_t2[95],s_t2[95]);
fa fau_1_96(b_i_s[96],s_t[96],c_t[95],c_t2[96],s_t2[96]);
fa fau_1_97(b_i_s[97],s_t[97],c_t[96],c_t2[97],s_t2[97]);
fa fau_1_98(b_i_s[98],s_t[98],c_t[97],c_t2[98],s_t2[98]);
fa fau_1_99(b_i_s[99],s_t[99],c_t[98],c_t2[99],s_t2[99]);
fa fau_1_100(b_i_s[100],s_t[100],c_t[99],c_t2[100],s_t2[100]);
fa fau_1_101(b_i_s[101],s_t[101],c_t[100],c_t2[101],s_t2[101]);
fa fau_1_102(b_i_s[102],s_t[102],c_t[101],c_t2[102],s_t2[102]);
fa fau_1_103(b_i_s[103],s_t[103],c_t[102],c_t2[103],s_t2[103]);
fa fau_1_104(b_i_s[104],s_t[104],c_t[103],c_t2[104],s_t2[104]);
fa fau_1_105(b_i_s[105],s_t[105],c_t[104],c_t2[105],s_t2[105]);
fa fau_1_106(b_i_s[106],s_t[106],c_t[105],c_t2[106],s_t2[106]);
fa fau_1_107(b_i_s[107],s_t[107],c_t[106],c_t2[107],s_t2[107]);
fa fau_1_108(b_i_s[108],s_t[108],c_t[107],c_t2[108],s_t2[108]);
fa fau_1_109(b_i_s[109],s_t[109],c_t[108],c_t2[109],s_t2[109]);
fa fau_1_110(b_i_s[110],s_t[110],c_t[109],c_t2[110],s_t2[110]);
fa fau_1_111(b_i_s[111],s_t[111],c_t[110],c_t2[111],s_t2[111]);
fa fau_1_112(b_i_s[112],s_t[112],c_t[111],c_t2[112],s_t2[112]);
fa fau_1_113(b_i_s[113],s_t[113],c_t[112],c_t2[113],s_t2[113]);
fa fau_1_114(b_i_s[114],s_t[114],c_t[113],c_t2[114],s_t2[114]);
fa fau_1_115(b_i_s[115],s_t[115],c_t[114],c_t2[115],s_t2[115]);
fa fau_1_116(b_i_s[116],s_t[116],c_t[115],c_t2[116],s_t2[116]);
fa fau_1_117(b_i_s[117],s_t[117],c_t[116],c_t2[117],s_t2[117]);
fa fau_1_118(b_i_s[118],s_t[118],c_t[117],c_t2[118],s_t2[118]);
fa fau_1_119(b_i_s[119],s_t[119],c_t[118],c_t2[119],s_t2[119]);
fa fau_1_120(b_i_s[120],s_t[120],c_t[119],c_t2[120],s_t2[120]);
fa fau_1_121(b_i_s[121],s_t[121],c_t[120],c_t2[121],s_t2[121]);
fa fau_1_122(b_i_s[122],s_t[122],c_t[121],c_t2[122],s_t2[122]);
fa fau_1_123(b_i_s[123],s_t[123],c_t[122],c_t2[123],s_t2[123]);
fa fau_1_124(b_i_s[124],s_t[124],c_t[123],c_t2[124],s_t2[124]);
fa fau_1_125(b_i_s[125],s_t[125],c_t[124],c_t2[125],s_t2[125]);
fa fau_1_126(b_i_s[126],s_t[126],c_t[125],c_t2[126],s_t2[126]);
fa fau_1_127(b_i_s[127],s_t[127],c_t[126],c_t2[127],s_t2[127]);
fa fau_1_128(b_i_s[128],s_t[128],c_t[127],c_t2[128],s_t2[128]);
fa fau_1_129(b_i_s[129],s_t[129],c_t[128],c_t2[129],s_t2[129]);
fa fau_1_130(b_i_s[130],s_t[130],c_t[129],c_t2[130],s_t2[130]);
fa fau_1_131(b_i_s[131],s_t[131],c_t[130],c_t2[131],s_t2[131]);
fa fau_1_132(b_i_s[132],s_t[132],c_t[131],c_t2[132],s_t2[132]);
fa fau_1_133(b_i_s[133],s_t[133],c_t[132],c_t2[133],s_t2[133]);
fa fau_1_134(b_i_s[134],s_t[134],c_t[133],c_t2[134],s_t2[134]);
fa fau_1_135(b_i_s[135],s_t[135],c_t[134],c_t2[135],s_t2[135]);
fa fau_1_136(b_i_s[136],s_t[136],c_t[135],c_t2[136],s_t2[136]);
fa fau_1_137(b_i_s[137],s_t[137],c_t[136],c_t2[137],s_t2[137]);
fa fau_1_138(b_i_s[138],s_t[138],c_t[137],c_t2[138],s_t2[138]);
fa fau_1_139(b_i_s[139],s_t[139],c_t[138],c_t2[139],s_t2[139]);
fa fau_1_140(b_i_s[140],s_t[140],c_t[139],c_t2[140],s_t2[140]);
fa fau_1_141(b_i_s[141],s_t[141],c_t[140],c_t2[141],s_t2[141]);
fa fau_1_142(b_i_s[142],s_t[142],c_t[141],c_t2[142],s_t2[142]);
fa fau_1_143(b_i_s[143],s_t[143],c_t[142],c_t2[143],s_t2[143]);
fa fau_1_144(b_i_s[144],s_t[144],c_t[143],c_t2[144],s_t2[144]);
fa fau_1_145(b_i_s[145],s_t[145],c_t[144],c_t2[145],s_t2[145]);
fa fau_1_146(b_i_s[146],s_t[146],c_t[145],c_t2[146],s_t2[146]);
fa fau_1_147(b_i_s[147],s_t[147],c_t[146],c_t2[147],s_t2[147]);
fa fau_1_148(b_i_s[148],s_t[148],c_t[147],c_t2[148],s_t2[148]);
fa fau_1_149(b_i_s[149],s_t[149],c_t[148],c_t2[149],s_t2[149]);
fa fau_1_150(b_i_s[150],s_t[150],c_t[149],c_t2[150],s_t2[150]);
fa fau_1_151(b_i_s[151],s_t[151],c_t[150],c_t2[151],s_t2[151]);
fa fau_1_152(b_i_s[152],s_t[152],c_t[151],c_t2[152],s_t2[152]);
fa fau_1_153(b_i_s[153],s_t[153],c_t[152],c_t2[153],s_t2[153]);
fa fau_1_154(b_i_s[154],s_t[154],c_t[153],c_t2[154],s_t2[154]);
fa fau_1_155(b_i_s[155],s_t[155],c_t[154],c_t2[155],s_t2[155]);
fa fau_1_156(b_i_s[156],s_t[156],c_t[155],c_t2[156],s_t2[156]);
fa fau_1_157(b_i_s[157],s_t[157],c_t[156],c_t2[157],s_t2[157]);
fa fau_1_158(b_i_s[158],s_t[158],c_t[157],c_t2[158],s_t2[158]);
fa fau_1_159(b_i_s[159],s_t[159],c_t[158],c_t2[159],s_t2[159]);
fa fau_1_160(b_i_s[160],s_t[160],c_t[159],c_t2[160],s_t2[160]);
fa fau_1_161(b_i_s[161],s_t[161],c_t[160],c_t2[161],s_t2[161]);
fa fau_1_162(b_i_s[162],s_t[162],c_t[161],c_t2[162],s_t2[162]);
fa fau_1_163(b_i_s[163],s_t[163],c_t[162],c_t2[163],s_t2[163]);
fa fau_1_164(b_i_s[164],s_t[164],c_t[163],c_t2[164],s_t2[164]);
fa fau_1_165(b_i_s[165],s_t[165],c_t[164],c_t2[165],s_t2[165]);
fa fau_1_166(b_i_s[166],s_t[166],c_t[165],c_t2[166],s_t2[166]);
fa fau_1_167(b_i_s[167],s_t[167],c_t[166],c_t2[167],s_t2[167]);
fa fau_1_168(b_i_s[168],s_t[168],c_t[167],c_t2[168],s_t2[168]);
fa fau_1_169(b_i_s[169],s_t[169],c_t[168],c_t2[169],s_t2[169]);
fa fau_1_170(b_i_s[170],s_t[170],c_t[169],c_t2[170],s_t2[170]);
fa fau_1_171(b_i_s[171],s_t[171],c_t[170],c_t2[171],s_t2[171]);
fa fau_1_172(b_i_s[172],s_t[172],c_t[171],c_t2[172],s_t2[172]);
fa fau_1_173(b_i_s[173],s_t[173],c_t[172],c_t2[173],s_t2[173]);
fa fau_1_174(b_i_s[174],s_t[174],c_t[173],c_t2[174],s_t2[174]);
fa fau_1_175(b_i_s[175],s_t[175],c_t[174],c_t2[175],s_t2[175]);
fa fau_1_176(b_i_s[176],s_t[176],c_t[175],c_t2[176],s_t2[176]);
fa fau_1_177(b_i_s[177],s_t[177],c_t[176],c_t2[177],s_t2[177]);
fa fau_1_178(b_i_s[178],s_t[178],c_t[177],c_t2[178],s_t2[178]);
fa fau_1_179(b_i_s[179],s_t[179],c_t[178],c_t2[179],s_t2[179]);
fa fau_1_180(b_i_s[180],s_t[180],c_t[179],c_t2[180],s_t2[180]);
fa fau_1_181(b_i_s[181],s_t[181],c_t[180],c_t2[181],s_t2[181]);
fa fau_1_182(b_i_s[182],s_t[182],c_t[181],c_t2[182],s_t2[182]);
fa fau_1_183(b_i_s[183],s_t[183],c_t[182],c_t2[183],s_t2[183]);
fa fau_1_184(b_i_s[184],s_t[184],c_t[183],c_t2[184],s_t2[184]);
fa fau_1_185(b_i_s[185],s_t[185],c_t[184],c_t2[185],s_t2[185]);
fa fau_1_186(b_i_s[186],s_t[186],c_t[185],c_t2[186],s_t2[186]);
fa fau_1_187(b_i_s[187],s_t[187],c_t[186],c_t2[187],s_t2[187]);
fa fau_1_188(b_i_s[188],s_t[188],c_t[187],c_t2[188],s_t2[188]);
fa fau_1_189(b_i_s[189],s_t[189],c_t[188],c_t2[189],s_t2[189]);
fa fau_1_190(b_i_s[190],s_t[190],c_t[189],c_t2[190],s_t2[190]);
fa fau_1_191(b_i_s[191],s_t[191],c_t[190],c_t2[191],s_t2[191]);
fa fau_1_192(b_i_s[192],s_t[192],c_t[191],c_t2[192],s_t2[192]);
fa fau_1_193(b_i_s[193],s_t[193],c_t[192],c_t2[193],s_t2[193]);
fa fau_1_194(b_i_s[194],s_t[194],c_t[193],c_t2[194],s_t2[194]);
fa fau_1_195(b_i_s[195],s_t[195],c_t[194],c_t2[195],s_t2[195]);
fa fau_1_196(b_i_s[196],s_t[196],c_t[195],c_t2[196],s_t2[196]);
fa fau_1_197(b_i_s[197],s_t[197],c_t[196],c_t2[197],s_t2[197]);
fa fau_1_198(b_i_s[198],s_t[198],c_t[197],c_t2[198],s_t2[198]);
fa fau_1_199(b_i_s[199],s_t[199],c_t[198],c_t2[199],s_t2[199]);
fa fau_1_200(b_i_s[200],s_t[200],c_t[199],c_t2[200],s_t2[200]);
fa fau_1_201(b_i_s[201],s_t[201],c_t[200],c_t2[201],s_t2[201]);
fa fau_1_202(b_i_s[202],s_t[202],c_t[201],c_t2[202],s_t2[202]);
fa fau_1_203(b_i_s[203],s_t[203],c_t[202],c_t2[203],s_t2[203]);
fa fau_1_204(b_i_s[204],s_t[204],c_t[203],c_t2[204],s_t2[204]);
fa fau_1_205(b_i_s[205],s_t[205],c_t[204],c_t2[205],s_t2[205]);
fa fau_1_206(b_i_s[206],s_t[206],c_t[205],c_t2[206],s_t2[206]);
fa fau_1_207(b_i_s[207],s_t[207],c_t[206],c_t2[207],s_t2[207]);
fa fau_1_208(b_i_s[208],s_t[208],c_t[207],c_t2[208],s_t2[208]);
fa fau_1_209(b_i_s[209],s_t[209],c_t[208],c_t2[209],s_t2[209]);
fa fau_1_210(b_i_s[210],s_t[210],c_t[209],c_t2[210],s_t2[210]);
fa fau_1_211(b_i_s[211],s_t[211],c_t[210],c_t2[211],s_t2[211]);
fa fau_1_212(b_i_s[212],s_t[212],c_t[211],c_t2[212],s_t2[212]);
fa fau_1_213(b_i_s[213],s_t[213],c_t[212],c_t2[213],s_t2[213]);
fa fau_1_214(b_i_s[214],s_t[214],c_t[213],c_t2[214],s_t2[214]);
fa fau_1_215(b_i_s[215],s_t[215],c_t[214],c_t2[215],s_t2[215]);
fa fau_1_216(b_i_s[216],s_t[216],c_t[215],c_t2[216],s_t2[216]);
fa fau_1_217(b_i_s[217],s_t[217],c_t[216],c_t2[217],s_t2[217]);
fa fau_1_218(b_i_s[218],s_t[218],c_t[217],c_t2[218],s_t2[218]);
fa fau_1_219(b_i_s[219],s_t[219],c_t[218],c_t2[219],s_t2[219]);
fa fau_1_220(b_i_s[220],s_t[220],c_t[219],c_t2[220],s_t2[220]);
fa fau_1_221(b_i_s[221],s_t[221],c_t[220],c_t2[221],s_t2[221]);
fa fau_1_222(b_i_s[222],s_t[222],c_t[221],c_t2[222],s_t2[222]);
fa fau_1_223(b_i_s[223],s_t[223],c_t[222],c_t2[223],s_t2[223]);
fa fau_1_224(b_i_s[224],s_t[224],c_t[223],c_t2[224],s_t2[224]);
fa fau_1_225(b_i_s[225],s_t[225],c_t[224],c_t2[225],s_t2[225]);
fa fau_1_226(b_i_s[226],s_t[226],c_t[225],c_t2[226],s_t2[226]);
fa fau_1_227(b_i_s[227],s_t[227],c_t[226],c_t2[227],s_t2[227]);
fa fau_1_228(b_i_s[228],s_t[228],c_t[227],c_t2[228],s_t2[228]);
fa fau_1_229(b_i_s[229],s_t[229],c_t[228],c_t2[229],s_t2[229]);
fa fau_1_230(b_i_s[230],s_t[230],c_t[229],c_t2[230],s_t2[230]);
fa fau_1_231(b_i_s[231],s_t[231],c_t[230],c_t2[231],s_t2[231]);
fa fau_1_232(b_i_s[232],s_t[232],c_t[231],c_t2[232],s_t2[232]);
fa fau_1_233(b_i_s[233],s_t[233],c_t[232],c_t2[233],s_t2[233]);
fa fau_1_234(b_i_s[234],s_t[234],c_t[233],c_t2[234],s_t2[234]);
fa fau_1_235(b_i_s[235],s_t[235],c_t[234],c_t2[235],s_t2[235]);
fa fau_1_236(b_i_s[236],s_t[236],c_t[235],c_t2[236],s_t2[236]);
fa fau_1_237(b_i_s[237],s_t[237],c_t[236],c_t2[237],s_t2[237]);
fa fau_1_238(b_i_s[238],s_t[238],c_t[237],c_t2[238],s_t2[238]);
fa fau_1_239(b_i_s[239],s_t[239],c_t[238],c_t2[239],s_t2[239]);
fa fau_1_240(b_i_s[240],s_t[240],c_t[239],c_t2[240],s_t2[240]);
fa fau_1_241(b_i_s[241],s_t[241],c_t[240],c_t2[241],s_t2[241]);
fa fau_1_242(b_i_s[242],s_t[242],c_t[241],c_t2[242],s_t2[242]);
fa fau_1_243(b_i_s[243],s_t[243],c_t[242],c_t2[243],s_t2[243]);
fa fau_1_244(b_i_s[244],s_t[244],c_t[243],c_t2[244],s_t2[244]);
fa fau_1_245(b_i_s[245],s_t[245],c_t[244],c_t2[245],s_t2[245]);
fa fau_1_246(b_i_s[246],s_t[246],c_t[245],c_t2[246],s_t2[246]);
fa fau_1_247(b_i_s[247],s_t[247],c_t[246],c_t2[247],s_t2[247]);
fa fau_1_248(b_i_s[248],s_t[248],c_t[247],c_t2[248],s_t2[248]);
fa fau_1_249(b_i_s[249],s_t[249],c_t[248],c_t2[249],s_t2[249]);
fa fau_1_250(b_i_s[250],s_t[250],c_t[249],c_t2[250],s_t2[250]);
fa fau_1_251(b_i_s[251],s_t[251],c_t[250],c_t2[251],s_t2[251]);
fa fau_1_252(b_i_s[252],s_t[252],c_t[251],c_t2[252],s_t2[252]);
fa fau_1_253(b_i_s[253],s_t[253],c_t[252],c_t2[253],s_t2[253]);
fa fau_1_254(b_i_s[254],s_t[254],c_t[253],c_t2[254],s_t2[254]);
fa fau_1_255(b_i_s[255],s_t[255],c_t[254],c_t2[255],s_t2[255]);
fa fau_1_256(b_i_s[256],s_t[256],c_t[255],c_t2[256],s_t2[256]);
fa fau_1_257(b_i_s[257],s_t[257],c_t[256],c_t2[257],s_t2[257]);
fa fau_1_258(b_i_s[258],s_t[258],c_t[257],c_t2[258],s_t2[258]);
fa fau_1_259(b_i_s[259],s_t[259],c_t[258],c_t2[259],s_t2[259]);
fa fau_1_260(b_i_s[260],s_t[260],c_t[259],c_t2[260],s_t2[260]);
fa fau_1_261(b_i_s[261],s_t[261],c_t[260],c_t2[261],s_t2[261]);
fa fau_1_262(b_i_s[262],s_t[262],c_t[261],c_t2[262],s_t2[262]);
fa fau_1_263(b_i_s[263],s_t[263],c_t[262],c_t2[263],s_t2[263]);
fa fau_1_264(b_i_s[264],s_t[264],c_t[263],c_t2[264],s_t2[264]);
fa fau_1_265(b_i_s[265],s_t[265],c_t[264],c_t2[265],s_t2[265]);
fa fau_1_266(b_i_s[266],s_t[266],c_t[265],c_t2[266],s_t2[266]);
fa fau_1_267(b_i_s[267],s_t[267],c_t[266],c_t2[267],s_t2[267]);
fa fau_1_268(b_i_s[268],s_t[268],c_t[267],c_t2[268],s_t2[268]);
fa fau_1_269(b_i_s[269],s_t[269],c_t[268],c_t2[269],s_t2[269]);
fa fau_1_270(b_i_s[270],s_t[270],c_t[269],c_t2[270],s_t2[270]);
fa fau_1_271(b_i_s[271],s_t[271],c_t[270],c_t2[271],s_t2[271]);
fa fau_1_272(b_i_s[272],s_t[272],c_t[271],c_t2[272],s_t2[272]);
fa fau_1_273(b_i_s[273],s_t[273],c_t[272],c_t2[273],s_t2[273]);
fa fau_1_274(b_i_s[274],s_t[274],c_t[273],c_t2[274],s_t2[274]);
fa fau_1_275(b_i_s[275],s_t[275],c_t[274],c_t2[275],s_t2[275]);
fa fau_1_276(b_i_s[276],s_t[276],c_t[275],c_t2[276],s_t2[276]);
fa fau_1_277(b_i_s[277],s_t[277],c_t[276],c_t2[277],s_t2[277]);
fa fau_1_278(b_i_s[278],s_t[278],c_t[277],c_t2[278],s_t2[278]);
fa fau_1_279(b_i_s[279],s_t[279],c_t[278],c_t2[279],s_t2[279]);
fa fau_1_280(b_i_s[280],s_t[280],c_t[279],c_t2[280],s_t2[280]);
fa fau_1_281(b_i_s[281],s_t[281],c_t[280],c_t2[281],s_t2[281]);
fa fau_1_282(b_i_s[282],s_t[282],c_t[281],c_t2[282],s_t2[282]);
fa fau_1_283(b_i_s[283],s_t[283],c_t[282],c_t2[283],s_t2[283]);
fa fau_1_284(b_i_s[284],s_t[284],c_t[283],c_t2[284],s_t2[284]);
fa fau_1_285(b_i_s[285],s_t[285],c_t[284],c_t2[285],s_t2[285]);
fa fau_1_286(b_i_s[286],s_t[286],c_t[285],c_t2[286],s_t2[286]);
fa fau_1_287(b_i_s[287],s_t[287],c_t[286],c_t2[287],s_t2[287]);
fa fau_1_288(b_i_s[288],s_t[288],c_t[287],c_t2[288],s_t2[288]);
fa fau_1_289(b_i_s[289],s_t[289],c_t[288],c_t2[289],s_t2[289]);
fa fau_1_290(b_i_s[290],s_t[290],c_t[289],c_t2[290],s_t2[290]);
fa fau_1_291(b_i_s[291],s_t[291],c_t[290],c_t2[291],s_t2[291]);
fa fau_1_292(b_i_s[292],s_t[292],c_t[291],c_t2[292],s_t2[292]);
fa fau_1_293(b_i_s[293],s_t[293],c_t[292],c_t2[293],s_t2[293]);
fa fau_1_294(b_i_s[294],s_t[294],c_t[293],c_t2[294],s_t2[294]);
fa fau_1_295(b_i_s[295],s_t[295],c_t[294],c_t2[295],s_t2[295]);
fa fau_1_296(b_i_s[296],s_t[296],c_t[295],c_t2[296],s_t2[296]);
fa fau_1_297(b_i_s[297],s_t[297],c_t[296],c_t2[297],s_t2[297]);
fa fau_1_298(b_i_s[298],s_t[298],c_t[297],c_t2[298],s_t2[298]);
fa fau_1_299(b_i_s[299],s_t[299],c_t[298],c_t2[299],s_t2[299]);
fa fau_1_300(b_i_s[300],s_t[300],c_t[299],c_t2[300],s_t2[300]);
fa fau_1_301(b_i_s[301],s_t[301],c_t[300],c_t2[301],s_t2[301]);
fa fau_1_302(b_i_s[302],s_t[302],c_t[301],c_t2[302],s_t2[302]);
fa fau_1_303(b_i_s[303],s_t[303],c_t[302],c_t2[303],s_t2[303]);
fa fau_1_304(b_i_s[304],s_t[304],c_t[303],c_t2[304],s_t2[304]);
fa fau_1_305(b_i_s[305],s_t[305],c_t[304],c_t2[305],s_t2[305]);
fa fau_1_306(b_i_s[306],s_t[306],c_t[305],c_t2[306],s_t2[306]);
fa fau_1_307(b_i_s[307],s_t[307],c_t[306],c_t2[307],s_t2[307]);
fa fau_1_308(b_i_s[308],s_t[308],c_t[307],c_t2[308],s_t2[308]);
fa fau_1_309(b_i_s[309],s_t[309],c_t[308],c_t2[309],s_t2[309]);
fa fau_1_310(b_i_s[310],s_t[310],c_t[309],c_t2[310],s_t2[310]);
fa fau_1_311(b_i_s[311],s_t[311],c_t[310],c_t2[311],s_t2[311]);
fa fau_1_312(b_i_s[312],s_t[312],c_t[311],c_t2[312],s_t2[312]);
fa fau_1_313(b_i_s[313],s_t[313],c_t[312],c_t2[313],s_t2[313]);
fa fau_1_314(b_i_s[314],s_t[314],c_t[313],c_t2[314],s_t2[314]);
fa fau_1_315(b_i_s[315],s_t[315],c_t[314],c_t2[315],s_t2[315]);
fa fau_1_316(b_i_s[316],s_t[316],c_t[315],c_t2[316],s_t2[316]);
fa fau_1_317(b_i_s[317],s_t[317],c_t[316],c_t2[317],s_t2[317]);
fa fau_1_318(b_i_s[318],s_t[318],c_t[317],c_t2[318],s_t2[318]);
fa fau_1_319(b_i_s[319],s_t[319],c_t[318],c_t2[319],s_t2[319]);
fa fau_1_320(b_i_s[320],s_t[320],c_t[319],c_t2[320],s_t2[320]);
fa fau_1_321(b_i_s[321],s_t[321],c_t[320],c_t2[321],s_t2[321]);
fa fau_1_322(b_i_s[322],s_t[322],c_t[321],c_t2[322],s_t2[322]);
fa fau_1_323(b_i_s[323],s_t[323],c_t[322],c_t2[323],s_t2[323]);
fa fau_1_324(b_i_s[324],s_t[324],c_t[323],c_t2[324],s_t2[324]);
fa fau_1_325(b_i_s[325],s_t[325],c_t[324],c_t2[325],s_t2[325]);
fa fau_1_326(b_i_s[326],s_t[326],c_t[325],c_t2[326],s_t2[326]);
fa fau_1_327(b_i_s[327],s_t[327],c_t[326],c_t2[327],s_t2[327]);
fa fau_1_328(b_i_s[328],s_t[328],c_t[327],c_t2[328],s_t2[328]);
fa fau_1_329(b_i_s[329],s_t[329],c_t[328],c_t2[329],s_t2[329]);
fa fau_1_330(b_i_s[330],s_t[330],c_t[329],c_t2[330],s_t2[330]);
fa fau_1_331(b_i_s[331],s_t[331],c_t[330],c_t2[331],s_t2[331]);
fa fau_1_332(b_i_s[332],s_t[332],c_t[331],c_t2[332],s_t2[332]);
fa fau_1_333(b_i_s[333],s_t[333],c_t[332],c_t2[333],s_t2[333]);
fa fau_1_334(b_i_s[334],s_t[334],c_t[333],c_t2[334],s_t2[334]);
fa fau_1_335(b_i_s[335],s_t[335],c_t[334],c_t2[335],s_t2[335]);
fa fau_1_336(b_i_s[336],s_t[336],c_t[335],c_t2[336],s_t2[336]);
fa fau_1_337(b_i_s[337],s_t[337],c_t[336],c_t2[337],s_t2[337]);
fa fau_1_338(b_i_s[338],s_t[338],c_t[337],c_t2[338],s_t2[338]);
fa fau_1_339(b_i_s[339],s_t[339],c_t[338],c_t2[339],s_t2[339]);
fa fau_1_340(b_i_s[340],s_t[340],c_t[339],c_t2[340],s_t2[340]);
fa fau_1_341(b_i_s[341],s_t[341],c_t[340],c_t2[341],s_t2[341]);
fa fau_1_342(b_i_s[342],s_t[342],c_t[341],c_t2[342],s_t2[342]);
fa fau_1_343(b_i_s[343],s_t[343],c_t[342],c_t2[343],s_t2[343]);
fa fau_1_344(b_i_s[344],s_t[344],c_t[343],c_t2[344],s_t2[344]);
fa fau_1_345(b_i_s[345],s_t[345],c_t[344],c_t2[345],s_t2[345]);
fa fau_1_346(b_i_s[346],s_t[346],c_t[345],c_t2[346],s_t2[346]);
fa fau_1_347(b_i_s[347],s_t[347],c_t[346],c_t2[347],s_t2[347]);
fa fau_1_348(b_i_s[348],s_t[348],c_t[347],c_t2[348],s_t2[348]);
fa fau_1_349(b_i_s[349],s_t[349],c_t[348],c_t2[349],s_t2[349]);
fa fau_1_350(b_i_s[350],s_t[350],c_t[349],c_t2[350],s_t2[350]);
fa fau_1_351(b_i_s[351],s_t[351],c_t[350],c_t2[351],s_t2[351]);
fa fau_1_352(b_i_s[352],s_t[352],c_t[351],c_t2[352],s_t2[352]);
fa fau_1_353(b_i_s[353],s_t[353],c_t[352],c_t2[353],s_t2[353]);
fa fau_1_354(b_i_s[354],s_t[354],c_t[353],c_t2[354],s_t2[354]);
fa fau_1_355(b_i_s[355],s_t[355],c_t[354],c_t2[355],s_t2[355]);
fa fau_1_356(b_i_s[356],s_t[356],c_t[355],c_t2[356],s_t2[356]);
fa fau_1_357(b_i_s[357],s_t[357],c_t[356],c_t2[357],s_t2[357]);
fa fau_1_358(b_i_s[358],s_t[358],c_t[357],c_t2[358],s_t2[358]);
fa fau_1_359(b_i_s[359],s_t[359],c_t[358],c_t2[359],s_t2[359]);
fa fau_1_360(b_i_s[360],s_t[360],c_t[359],c_t2[360],s_t2[360]);
fa fau_1_361(b_i_s[361],s_t[361],c_t[360],c_t2[361],s_t2[361]);
fa fau_1_362(b_i_s[362],s_t[362],c_t[361],c_t2[362],s_t2[362]);
fa fau_1_363(b_i_s[363],s_t[363],c_t[362],c_t2[363],s_t2[363]);
fa fau_1_364(b_i_s[364],s_t[364],c_t[363],c_t2[364],s_t2[364]);
fa fau_1_365(b_i_s[365],s_t[365],c_t[364],c_t2[365],s_t2[365]);
fa fau_1_366(b_i_s[366],s_t[366],c_t[365],c_t2[366],s_t2[366]);
fa fau_1_367(b_i_s[367],s_t[367],c_t[366],c_t2[367],s_t2[367]);
fa fau_1_368(b_i_s[368],s_t[368],c_t[367],c_t2[368],s_t2[368]);
fa fau_1_369(b_i_s[369],s_t[369],c_t[368],c_t2[369],s_t2[369]);
fa fau_1_370(b_i_s[370],s_t[370],c_t[369],c_t2[370],s_t2[370]);
fa fau_1_371(b_i_s[371],s_t[371],c_t[370],c_t2[371],s_t2[371]);
fa fau_1_372(b_i_s[372],s_t[372],c_t[371],c_t2[372],s_t2[372]);
fa fau_1_373(b_i_s[373],s_t[373],c_t[372],c_t2[373],s_t2[373]);
fa fau_1_374(b_i_s[374],s_t[374],c_t[373],c_t2[374],s_t2[374]);
fa fau_1_375(b_i_s[375],s_t[375],c_t[374],c_t2[375],s_t2[375]);
fa fau_1_376(b_i_s[376],s_t[376],c_t[375],c_t2[376],s_t2[376]);
fa fau_1_377(b_i_s[377],s_t[377],c_t[376],c_t2[377],s_t2[377]);
fa fau_1_378(b_i_s[378],s_t[378],c_t[377],c_t2[378],s_t2[378]);
fa fau_1_379(b_i_s[379],s_t[379],c_t[378],c_t2[379],s_t2[379]);
fa fau_1_380(b_i_s[380],s_t[380],c_t[379],c_t2[380],s_t2[380]);
fa fau_1_381(b_i_s[381],s_t[381],c_t[380],c_t2[381],s_t2[381]);
fa fau_1_382(b_i_s[382],s_t[382],c_t[381],c_t2[382],s_t2[382]);
fa fau_1_383(b_i_s[383],s_t[383],c_t[382],c_t2[383],s_t2[383]);
fa fau_1_384(b_i_s[384],s_t[384],c_t[383],c_t2[384],s_t2[384]);
fa fau_1_385(b_i_s[385],s_t[385],c_t[384],c_t2[385],s_t2[385]);
fa fau_1_386(b_i_s[386],s_t[386],c_t[385],c_t2[386],s_t2[386]);
fa fau_1_387(b_i_s[387],s_t[387],c_t[386],c_t2[387],s_t2[387]);
fa fau_1_388(b_i_s[388],s_t[388],c_t[387],c_t2[388],s_t2[388]);
fa fau_1_389(b_i_s[389],s_t[389],c_t[388],c_t2[389],s_t2[389]);
fa fau_1_390(b_i_s[390],s_t[390],c_t[389],c_t2[390],s_t2[390]);
fa fau_1_391(b_i_s[391],s_t[391],c_t[390],c_t2[391],s_t2[391]);
fa fau_1_392(b_i_s[392],s_t[392],c_t[391],c_t2[392],s_t2[392]);
fa fau_1_393(b_i_s[393],s_t[393],c_t[392],c_t2[393],s_t2[393]);
fa fau_1_394(b_i_s[394],s_t[394],c_t[393],c_t2[394],s_t2[394]);
fa fau_1_395(b_i_s[395],s_t[395],c_t[394],c_t2[395],s_t2[395]);
fa fau_1_396(b_i_s[396],s_t[396],c_t[395],c_t2[396],s_t2[396]);
fa fau_1_397(b_i_s[397],s_t[397],c_t[396],c_t2[397],s_t2[397]);
fa fau_1_398(b_i_s[398],s_t[398],c_t[397],c_t2[398],s_t2[398]);
fa fau_1_399(b_i_s[399],s_t[399],c_t[398],c_t2[399],s_t2[399]);
fa fau_1_400(b_i_s[400],s_t[400],c_t[399],c_t2[400],s_t2[400]);
fa fau_1_401(b_i_s[401],s_t[401],c_t[400],c_t2[401],s_t2[401]);
fa fau_1_402(b_i_s[402],s_t[402],c_t[401],c_t2[402],s_t2[402]);
fa fau_1_403(b_i_s[403],s_t[403],c_t[402],c_t2[403],s_t2[403]);
fa fau_1_404(b_i_s[404],s_t[404],c_t[403],c_t2[404],s_t2[404]);
fa fau_1_405(b_i_s[405],s_t[405],c_t[404],c_t2[405],s_t2[405]);
fa fau_1_406(b_i_s[406],s_t[406],c_t[405],c_t2[406],s_t2[406]);
fa fau_1_407(b_i_s[407],s_t[407],c_t[406],c_t2[407],s_t2[407]);
fa fau_1_408(b_i_s[408],s_t[408],c_t[407],c_t2[408],s_t2[408]);
fa fau_1_409(b_i_s[409],s_t[409],c_t[408],c_t2[409],s_t2[409]);
fa fau_1_410(b_i_s[410],s_t[410],c_t[409],c_t2[410],s_t2[410]);
fa fau_1_411(b_i_s[411],s_t[411],c_t[410],c_t2[411],s_t2[411]);
fa fau_1_412(b_i_s[412],s_t[412],c_t[411],c_t2[412],s_t2[412]);
fa fau_1_413(b_i_s[413],s_t[413],c_t[412],c_t2[413],s_t2[413]);
fa fau_1_414(b_i_s[414],s_t[414],c_t[413],c_t2[414],s_t2[414]);
fa fau_1_415(b_i_s[415],s_t[415],c_t[414],c_t2[415],s_t2[415]);
fa fau_1_416(b_i_s[416],s_t[416],c_t[415],c_t2[416],s_t2[416]);
fa fau_1_417(b_i_s[417],s_t[417],c_t[416],c_t2[417],s_t2[417]);
fa fau_1_418(b_i_s[418],s_t[418],c_t[417],c_t2[418],s_t2[418]);
fa fau_1_419(b_i_s[419],s_t[419],c_t[418],c_t2[419],s_t2[419]);
fa fau_1_420(b_i_s[420],s_t[420],c_t[419],c_t2[420],s_t2[420]);
fa fau_1_421(b_i_s[421],s_t[421],c_t[420],c_t2[421],s_t2[421]);
fa fau_1_422(b_i_s[422],s_t[422],c_t[421],c_t2[422],s_t2[422]);
fa fau_1_423(b_i_s[423],s_t[423],c_t[422],c_t2[423],s_t2[423]);
fa fau_1_424(b_i_s[424],s_t[424],c_t[423],c_t2[424],s_t2[424]);
fa fau_1_425(b_i_s[425],s_t[425],c_t[424],c_t2[425],s_t2[425]);
fa fau_1_426(b_i_s[426],s_t[426],c_t[425],c_t2[426],s_t2[426]);
fa fau_1_427(b_i_s[427],s_t[427],c_t[426],c_t2[427],s_t2[427]);
fa fau_1_428(b_i_s[428],s_t[428],c_t[427],c_t2[428],s_t2[428]);
fa fau_1_429(b_i_s[429],s_t[429],c_t[428],c_t2[429],s_t2[429]);
fa fau_1_430(b_i_s[430],s_t[430],c_t[429],c_t2[430],s_t2[430]);
fa fau_1_431(b_i_s[431],s_t[431],c_t[430],c_t2[431],s_t2[431]);
fa fau_1_432(b_i_s[432],s_t[432],c_t[431],c_t2[432],s_t2[432]);
fa fau_1_433(b_i_s[433],s_t[433],c_t[432],c_t2[433],s_t2[433]);
fa fau_1_434(b_i_s[434],s_t[434],c_t[433],c_t2[434],s_t2[434]);
fa fau_1_435(b_i_s[435],s_t[435],c_t[434],c_t2[435],s_t2[435]);
fa fau_1_436(b_i_s[436],s_t[436],c_t[435],c_t2[436],s_t2[436]);
fa fau_1_437(b_i_s[437],s_t[437],c_t[436],c_t2[437],s_t2[437]);
fa fau_1_438(b_i_s[438],s_t[438],c_t[437],c_t2[438],s_t2[438]);
fa fau_1_439(b_i_s[439],s_t[439],c_t[438],c_t2[439],s_t2[439]);
fa fau_1_440(b_i_s[440],s_t[440],c_t[439],c_t2[440],s_t2[440]);
fa fau_1_441(b_i_s[441],s_t[441],c_t[440],c_t2[441],s_t2[441]);
fa fau_1_442(b_i_s[442],s_t[442],c_t[441],c_t2[442],s_t2[442]);
fa fau_1_443(b_i_s[443],s_t[443],c_t[442],c_t2[443],s_t2[443]);
fa fau_1_444(b_i_s[444],s_t[444],c_t[443],c_t2[444],s_t2[444]);
fa fau_1_445(b_i_s[445],s_t[445],c_t[444],c_t2[445],s_t2[445]);
fa fau_1_446(b_i_s[446],s_t[446],c_t[445],c_t2[446],s_t2[446]);
fa fau_1_447(b_i_s[447],s_t[447],c_t[446],c_t2[447],s_t2[447]);
fa fau_1_448(b_i_s[448],s_t[448],c_t[447],c_t2[448],s_t2[448]);
fa fau_1_449(b_i_s[449],s_t[449],c_t[448],c_t2[449],s_t2[449]);
fa fau_1_450(b_i_s[450],s_t[450],c_t[449],c_t2[450],s_t2[450]);
fa fau_1_451(b_i_s[451],s_t[451],c_t[450],c_t2[451],s_t2[451]);
fa fau_1_452(b_i_s[452],s_t[452],c_t[451],c_t2[452],s_t2[452]);
fa fau_1_453(b_i_s[453],s_t[453],c_t[452],c_t2[453],s_t2[453]);
fa fau_1_454(b_i_s[454],s_t[454],c_t[453],c_t2[454],s_t2[454]);
fa fau_1_455(b_i_s[455],s_t[455],c_t[454],c_t2[455],s_t2[455]);
fa fau_1_456(b_i_s[456],s_t[456],c_t[455],c_t2[456],s_t2[456]);
fa fau_1_457(b_i_s[457],s_t[457],c_t[456],c_t2[457],s_t2[457]);
fa fau_1_458(b_i_s[458],s_t[458],c_t[457],c_t2[458],s_t2[458]);
fa fau_1_459(b_i_s[459],s_t[459],c_t[458],c_t2[459],s_t2[459]);
fa fau_1_460(b_i_s[460],s_t[460],c_t[459],c_t2[460],s_t2[460]);
fa fau_1_461(b_i_s[461],s_t[461],c_t[460],c_t2[461],s_t2[461]);
fa fau_1_462(b_i_s[462],s_t[462],c_t[461],c_t2[462],s_t2[462]);
fa fau_1_463(b_i_s[463],s_t[463],c_t[462],c_t2[463],s_t2[463]);
fa fau_1_464(b_i_s[464],s_t[464],c_t[463],c_t2[464],s_t2[464]);
fa fau_1_465(b_i_s[465],s_t[465],c_t[464],c_t2[465],s_t2[465]);
fa fau_1_466(b_i_s[466],s_t[466],c_t[465],c_t2[466],s_t2[466]);
fa fau_1_467(b_i_s[467],s_t[467],c_t[466],c_t2[467],s_t2[467]);
fa fau_1_468(b_i_s[468],s_t[468],c_t[467],c_t2[468],s_t2[468]);
fa fau_1_469(b_i_s[469],s_t[469],c_t[468],c_t2[469],s_t2[469]);
fa fau_1_470(b_i_s[470],s_t[470],c_t[469],c_t2[470],s_t2[470]);
fa fau_1_471(b_i_s[471],s_t[471],c_t[470],c_t2[471],s_t2[471]);
fa fau_1_472(b_i_s[472],s_t[472],c_t[471],c_t2[472],s_t2[472]);
fa fau_1_473(b_i_s[473],s_t[473],c_t[472],c_t2[473],s_t2[473]);
fa fau_1_474(b_i_s[474],s_t[474],c_t[473],c_t2[474],s_t2[474]);
fa fau_1_475(b_i_s[475],s_t[475],c_t[474],c_t2[475],s_t2[475]);
fa fau_1_476(b_i_s[476],s_t[476],c_t[475],c_t2[476],s_t2[476]);
fa fau_1_477(b_i_s[477],s_t[477],c_t[476],c_t2[477],s_t2[477]);
fa fau_1_478(b_i_s[478],s_t[478],c_t[477],c_t2[478],s_t2[478]);
fa fau_1_479(b_i_s[479],s_t[479],c_t[478],c_t2[479],s_t2[479]);
fa fau_1_480(b_i_s[480],s_t[480],c_t[479],c_t2[480],s_t2[480]);
fa fau_1_481(b_i_s[481],s_t[481],c_t[480],c_t2[481],s_t2[481]);
fa fau_1_482(b_i_s[482],s_t[482],c_t[481],c_t2[482],s_t2[482]);
fa fau_1_483(b_i_s[483],s_t[483],c_t[482],c_t2[483],s_t2[483]);
fa fau_1_484(b_i_s[484],s_t[484],c_t[483],c_t2[484],s_t2[484]);
fa fau_1_485(b_i_s[485],s_t[485],c_t[484],c_t2[485],s_t2[485]);
fa fau_1_486(b_i_s[486],s_t[486],c_t[485],c_t2[486],s_t2[486]);
fa fau_1_487(b_i_s[487],s_t[487],c_t[486],c_t2[487],s_t2[487]);
fa fau_1_488(b_i_s[488],s_t[488],c_t[487],c_t2[488],s_t2[488]);
fa fau_1_489(b_i_s[489],s_t[489],c_t[488],c_t2[489],s_t2[489]);
fa fau_1_490(b_i_s[490],s_t[490],c_t[489],c_t2[490],s_t2[490]);
fa fau_1_491(b_i_s[491],s_t[491],c_t[490],c_t2[491],s_t2[491]);
fa fau_1_492(b_i_s[492],s_t[492],c_t[491],c_t2[492],s_t2[492]);
fa fau_1_493(b_i_s[493],s_t[493],c_t[492],c_t2[493],s_t2[493]);
fa fau_1_494(b_i_s[494],s_t[494],c_t[493],c_t2[494],s_t2[494]);
fa fau_1_495(b_i_s[495],s_t[495],c_t[494],c_t2[495],s_t2[495]);
fa fau_1_496(b_i_s[496],s_t[496],c_t[495],c_t2[496],s_t2[496]);
fa fau_1_497(b_i_s[497],s_t[497],c_t[496],c_t2[497],s_t2[497]);
fa fau_1_498(b_i_s[498],s_t[498],c_t[497],c_t2[498],s_t2[498]);
fa fau_1_499(b_i_s[499],s_t[499],c_t[498],c_t2[499],s_t2[499]);
fa fau_1_500(b_i_s[500],s_t[500],c_t[499],c_t2[500],s_t2[500]);
fa fau_1_501(b_i_s[501],s_t[501],c_t[500],c_t2[501],s_t2[501]);
fa fau_1_502(b_i_s[502],s_t[502],c_t[501],c_t2[502],s_t2[502]);
fa fau_1_503(b_i_s[503],s_t[503],c_t[502],c_t2[503],s_t2[503]);
fa fau_1_504(b_i_s[504],s_t[504],c_t[503],c_t2[504],s_t2[504]);
fa fau_1_505(b_i_s[505],s_t[505],c_t[504],c_t2[505],s_t2[505]);
fa fau_1_506(b_i_s[506],s_t[506],c_t[505],c_t2[506],s_t2[506]);
fa fau_1_507(b_i_s[507],s_t[507],c_t[506],c_t2[507],s_t2[507]);
fa fau_1_508(b_i_s[508],s_t[508],c_t[507],c_t2[508],s_t2[508]);
fa fau_1_509(b_i_s[509],s_t[509],c_t[508],c_t2[509],s_t2[509]);
fa fau_1_510(b_i_s[510],s_t[510],c_t[509],c_t2[510],s_t2[510]);
fa fau_1_511(b_i_s[511],s_t[511],c_t[510],c_t2[511],s_t2[511]);
fa fau_1_512(b_i_s[512],s_t[512],c_t[511],c_t2[512],s_t2[512]);
fa fau_1_513(b_i_s[513],s_t[513],c_t[512],c_t2[513],s_t2[513]);
fa fau_1_514(b_i_s[514],s_t[514],c_t[513],c_t2[514],s_t2[514]);
fa fau_1_515(b_i_s[515],s_t[515],c_t[514],c_t2[515],s_t2[515]);
fa fau_1_516(b_i_s[516],s_t[516],c_t[515],c_t2[516],s_t2[516]);
fa fau_1_517(b_i_s[517],s_t[517],c_t[516],c_t2[517],s_t2[517]);
fa fau_1_518(b_i_s[518],s_t[518],c_t[517],c_t2[518],s_t2[518]);
fa fau_1_519(b_i_s[519],s_t[519],c_t[518],c_t2[519],s_t2[519]);
fa fau_1_520(b_i_s[520],s_t[520],c_t[519],c_t2[520],s_t2[520]);
fa fau_1_521(b_i_s[521],s_t[521],c_t[520],c_t2[521],s_t2[521]);
fa fau_1_522(b_i_s[522],s_t[522],c_t[521],c_t2[522],s_t2[522]);
fa fau_1_523(b_i_s[523],s_t[523],c_t[522],c_t2[523],s_t2[523]);
fa fau_1_524(b_i_s[524],s_t[524],c_t[523],c_t2[524],s_t2[524]);
fa fau_1_525(b_i_s[525],s_t[525],c_t[524],c_t2[525],s_t2[525]);
fa fau_1_526(b_i_s[526],s_t[526],c_t[525],c_t2[526],s_t2[526]);
fa fau_1_527(b_i_s[527],s_t[527],c_t[526],c_t2[527],s_t2[527]);
fa fau_1_528(b_i_s[528],s_t[528],c_t[527],c_t2[528],s_t2[528]);
fa fau_1_529(b_i_s[529],s_t[529],c_t[528],c_t2[529],s_t2[529]);
fa fau_1_530(b_i_s[530],s_t[530],c_t[529],c_t2[530],s_t2[530]);
fa fau_1_531(b_i_s[531],s_t[531],c_t[530],c_t2[531],s_t2[531]);
fa fau_1_532(b_i_s[532],s_t[532],c_t[531],c_t2[532],s_t2[532]);
fa fau_1_533(b_i_s[533],s_t[533],c_t[532],c_t2[533],s_t2[533]);
fa fau_1_534(b_i_s[534],s_t[534],c_t[533],c_t2[534],s_t2[534]);
fa fau_1_535(b_i_s[535],s_t[535],c_t[534],c_t2[535],s_t2[535]);
fa fau_1_536(b_i_s[536],s_t[536],c_t[535],c_t2[536],s_t2[536]);
fa fau_1_537(b_i_s[537],s_t[537],c_t[536],c_t2[537],s_t2[537]);
fa fau_1_538(b_i_s[538],s_t[538],c_t[537],c_t2[538],s_t2[538]);
fa fau_1_539(b_i_s[539],s_t[539],c_t[538],c_t2[539],s_t2[539]);
fa fau_1_540(b_i_s[540],s_t[540],c_t[539],c_t2[540],s_t2[540]);
fa fau_1_541(b_i_s[541],s_t[541],c_t[540],c_t2[541],s_t2[541]);
fa fau_1_542(b_i_s[542],s_t[542],c_t[541],c_t2[542],s_t2[542]);
fa fau_1_543(b_i_s[543],s_t[543],c_t[542],c_t2[543],s_t2[543]);
fa fau_1_544(b_i_s[544],s_t[544],c_t[543],c_t2[544],s_t2[544]);
fa fau_1_545(b_i_s[545],s_t[545],c_t[544],c_t2[545],s_t2[545]);
fa fau_1_546(b_i_s[546],s_t[546],c_t[545],c_t2[546],s_t2[546]);
fa fau_1_547(b_i_s[547],s_t[547],c_t[546],c_t2[547],s_t2[547]);
fa fau_1_548(b_i_s[548],s_t[548],c_t[547],c_t2[548],s_t2[548]);
fa fau_1_549(b_i_s[549],s_t[549],c_t[548],c_t2[549],s_t2[549]);
fa fau_1_550(b_i_s[550],s_t[550],c_t[549],c_t2[550],s_t2[550]);
fa fau_1_551(b_i_s[551],s_t[551],c_t[550],c_t2[551],s_t2[551]);
fa fau_1_552(b_i_s[552],s_t[552],c_t[551],c_t2[552],s_t2[552]);
fa fau_1_553(b_i_s[553],s_t[553],c_t[552],c_t2[553],s_t2[553]);
fa fau_1_554(b_i_s[554],s_t[554],c_t[553],c_t2[554],s_t2[554]);
fa fau_1_555(b_i_s[555],s_t[555],c_t[554],c_t2[555],s_t2[555]);
fa fau_1_556(b_i_s[556],s_t[556],c_t[555],c_t2[556],s_t2[556]);
fa fau_1_557(b_i_s[557],s_t[557],c_t[556],c_t2[557],s_t2[557]);
fa fau_1_558(b_i_s[558],s_t[558],c_t[557],c_t2[558],s_t2[558]);
fa fau_1_559(b_i_s[559],s_t[559],c_t[558],c_t2[559],s_t2[559]);
fa fau_1_560(b_i_s[560],s_t[560],c_t[559],c_t2[560],s_t2[560]);
fa fau_1_561(b_i_s[561],s_t[561],c_t[560],c_t2[561],s_t2[561]);
fa fau_1_562(b_i_s[562],s_t[562],c_t[561],c_t2[562],s_t2[562]);
fa fau_1_563(b_i_s[563],s_t[563],c_t[562],c_t2[563],s_t2[563]);
fa fau_1_564(b_i_s[564],s_t[564],c_t[563],c_t2[564],s_t2[564]);
fa fau_1_565(b_i_s[565],s_t[565],c_t[564],c_t2[565],s_t2[565]);
fa fau_1_566(b_i_s[566],s_t[566],c_t[565],c_t2[566],s_t2[566]);
fa fau_1_567(b_i_s[567],s_t[567],c_t[566],c_t2[567],s_t2[567]);
fa fau_1_568(b_i_s[568],s_t[568],c_t[567],c_t2[568],s_t2[568]);
fa fau_1_569(b_i_s[569],s_t[569],c_t[568],c_t2[569],s_t2[569]);
fa fau_1_570(b_i_s[570],s_t[570],c_t[569],c_t2[570],s_t2[570]);
fa fau_1_571(b_i_s[571],s_t[571],c_t[570],c_t2[571],s_t2[571]);
fa fau_1_572(b_i_s[572],s_t[572],c_t[571],c_t2[572],s_t2[572]);
fa fau_1_573(b_i_s[573],s_t[573],c_t[572],c_t2[573],s_t2[573]);
fa fau_1_574(b_i_s[574],s_t[574],c_t[573],c_t2[574],s_t2[574]);
fa fau_1_575(b_i_s[575],s_t[575],c_t[574],c_t2[575],s_t2[575]);
fa fau_1_576(b_i_s[576],s_t[576],c_t[575],c_t2[576],s_t2[576]);
fa fau_1_577(b_i_s[577],s_t[577],c_t[576],c_t2[577],s_t2[577]);
fa fau_1_578(b_i_s[578],s_t[578],c_t[577],c_t2[578],s_t2[578]);
fa fau_1_579(b_i_s[579],s_t[579],c_t[578],c_t2[579],s_t2[579]);
fa fau_1_580(b_i_s[580],s_t[580],c_t[579],c_t2[580],s_t2[580]);
fa fau_1_581(b_i_s[581],s_t[581],c_t[580],c_t2[581],s_t2[581]);
fa fau_1_582(b_i_s[582],s_t[582],c_t[581],c_t2[582],s_t2[582]);
fa fau_1_583(b_i_s[583],s_t[583],c_t[582],c_t2[583],s_t2[583]);
fa fau_1_584(b_i_s[584],s_t[584],c_t[583],c_t2[584],s_t2[584]);
fa fau_1_585(b_i_s[585],s_t[585],c_t[584],c_t2[585],s_t2[585]);
fa fau_1_586(b_i_s[586],s_t[586],c_t[585],c_t2[586],s_t2[586]);
fa fau_1_587(b_i_s[587],s_t[587],c_t[586],c_t2[587],s_t2[587]);
fa fau_1_588(b_i_s[588],s_t[588],c_t[587],c_t2[588],s_t2[588]);
fa fau_1_589(b_i_s[589],s_t[589],c_t[588],c_t2[589],s_t2[589]);
fa fau_1_590(b_i_s[590],s_t[590],c_t[589],c_t2[590],s_t2[590]);
fa fau_1_591(b_i_s[591],s_t[591],c_t[590],c_t2[591],s_t2[591]);
fa fau_1_592(b_i_s[592],s_t[592],c_t[591],c_t2[592],s_t2[592]);
fa fau_1_593(b_i_s[593],s_t[593],c_t[592],c_t2[593],s_t2[593]);
fa fau_1_594(b_i_s[594],s_t[594],c_t[593],c_t2[594],s_t2[594]);
fa fau_1_595(b_i_s[595],s_t[595],c_t[594],c_t2[595],s_t2[595]);
fa fau_1_596(b_i_s[596],s_t[596],c_t[595],c_t2[596],s_t2[596]);
fa fau_1_597(b_i_s[597],s_t[597],c_t[596],c_t2[597],s_t2[597]);
fa fau_1_598(b_i_s[598],s_t[598],c_t[597],c_t2[598],s_t2[598]);
fa fau_1_599(b_i_s[599],s_t[599],c_t[598],c_t2[599],s_t2[599]);
fa fau_1_600(b_i_s[600],s_t[600],c_t[599],c_t2[600],s_t2[600]);
fa fau_1_601(b_i_s[601],s_t[601],c_t[600],c_t2[601],s_t2[601]);
fa fau_1_602(b_i_s[602],s_t[602],c_t[601],c_t2[602],s_t2[602]);
fa fau_1_603(b_i_s[603],s_t[603],c_t[602],c_t2[603],s_t2[603]);
fa fau_1_604(b_i_s[604],s_t[604],c_t[603],c_t2[604],s_t2[604]);
fa fau_1_605(b_i_s[605],s_t[605],c_t[604],c_t2[605],s_t2[605]);
fa fau_1_606(b_i_s[606],s_t[606],c_t[605],c_t2[606],s_t2[606]);
fa fau_1_607(b_i_s[607],s_t[607],c_t[606],c_t2[607],s_t2[607]);
fa fau_1_608(b_i_s[608],s_t[608],c_t[607],c_t2[608],s_t2[608]);
fa fau_1_609(b_i_s[609],s_t[609],c_t[608],c_t2[609],s_t2[609]);
fa fau_1_610(b_i_s[610],s_t[610],c_t[609],c_t2[610],s_t2[610]);
fa fau_1_611(b_i_s[611],s_t[611],c_t[610],c_t2[611],s_t2[611]);
fa fau_1_612(b_i_s[612],s_t[612],c_t[611],c_t2[612],s_t2[612]);
fa fau_1_613(b_i_s[613],s_t[613],c_t[612],c_t2[613],s_t2[613]);
fa fau_1_614(b_i_s[614],s_t[614],c_t[613],c_t2[614],s_t2[614]);
fa fau_1_615(b_i_s[615],s_t[615],c_t[614],c_t2[615],s_t2[615]);
fa fau_1_616(b_i_s[616],s_t[616],c_t[615],c_t2[616],s_t2[616]);
fa fau_1_617(b_i_s[617],s_t[617],c_t[616],c_t2[617],s_t2[617]);
fa fau_1_618(b_i_s[618],s_t[618],c_t[617],c_t2[618],s_t2[618]);
fa fau_1_619(b_i_s[619],s_t[619],c_t[618],c_t2[619],s_t2[619]);
fa fau_1_620(b_i_s[620],s_t[620],c_t[619],c_t2[620],s_t2[620]);
fa fau_1_621(b_i_s[621],s_t[621],c_t[620],c_t2[621],s_t2[621]);
fa fau_1_622(b_i_s[622],s_t[622],c_t[621],c_t2[622],s_t2[622]);
fa fau_1_623(b_i_s[623],s_t[623],c_t[622],c_t2[623],s_t2[623]);
fa fau_1_624(b_i_s[624],s_t[624],c_t[623],c_t2[624],s_t2[624]);
fa fau_1_625(b_i_s[625],s_t[625],c_t[624],c_t2[625],s_t2[625]);
fa fau_1_626(b_i_s[626],s_t[626],c_t[625],c_t2[626],s_t2[626]);
fa fau_1_627(b_i_s[627],s_t[627],c_t[626],c_t2[627],s_t2[627]);
fa fau_1_628(b_i_s[628],s_t[628],c_t[627],c_t2[628],s_t2[628]);
fa fau_1_629(b_i_s[629],s_t[629],c_t[628],c_t2[629],s_t2[629]);
fa fau_1_630(b_i_s[630],s_t[630],c_t[629],c_t2[630],s_t2[630]);
fa fau_1_631(b_i_s[631],s_t[631],c_t[630],c_t2[631],s_t2[631]);
fa fau_1_632(b_i_s[632],s_t[632],c_t[631],c_t2[632],s_t2[632]);
fa fau_1_633(b_i_s[633],s_t[633],c_t[632],c_t2[633],s_t2[633]);
fa fau_1_634(b_i_s[634],s_t[634],c_t[633],c_t2[634],s_t2[634]);
fa fau_1_635(b_i_s[635],s_t[635],c_t[634],c_t2[635],s_t2[635]);
fa fau_1_636(b_i_s[636],s_t[636],c_t[635],c_t2[636],s_t2[636]);
fa fau_1_637(b_i_s[637],s_t[637],c_t[636],c_t2[637],s_t2[637]);
fa fau_1_638(b_i_s[638],s_t[638],c_t[637],c_t2[638],s_t2[638]);
fa fau_1_639(b_i_s[639],s_t[639],c_t[638],c_t2[639],s_t2[639]);
fa fau_1_640(b_i_s[640],s_t[640],c_t[639],c_t2[640],s_t2[640]);
fa fau_1_641(b_i_s[641],s_t[641],c_t[640],c_t2[641],s_t2[641]);
fa fau_1_642(b_i_s[642],s_t[642],c_t[641],c_t2[642],s_t2[642]);
fa fau_1_643(b_i_s[643],s_t[643],c_t[642],c_t2[643],s_t2[643]);
fa fau_1_644(b_i_s[644],s_t[644],c_t[643],c_t2[644],s_t2[644]);
fa fau_1_645(b_i_s[645],s_t[645],c_t[644],c_t2[645],s_t2[645]);
fa fau_1_646(b_i_s[646],s_t[646],c_t[645],c_t2[646],s_t2[646]);
fa fau_1_647(b_i_s[647],s_t[647],c_t[646],c_t2[647],s_t2[647]);
fa fau_1_648(b_i_s[648],s_t[648],c_t[647],c_t2[648],s_t2[648]);
fa fau_1_649(b_i_s[649],s_t[649],c_t[648],c_t2[649],s_t2[649]);
fa fau_1_650(b_i_s[650],s_t[650],c_t[649],c_t2[650],s_t2[650]);
fa fau_1_651(b_i_s[651],s_t[651],c_t[650],c_t2[651],s_t2[651]);
fa fau_1_652(b_i_s[652],s_t[652],c_t[651],c_t2[652],s_t2[652]);
fa fau_1_653(b_i_s[653],s_t[653],c_t[652],c_t2[653],s_t2[653]);
fa fau_1_654(b_i_s[654],s_t[654],c_t[653],c_t2[654],s_t2[654]);
fa fau_1_655(b_i_s[655],s_t[655],c_t[654],c_t2[655],s_t2[655]);
fa fau_1_656(b_i_s[656],s_t[656],c_t[655],c_t2[656],s_t2[656]);
fa fau_1_657(b_i_s[657],s_t[657],c_t[656],c_t2[657],s_t2[657]);
fa fau_1_658(b_i_s[658],s_t[658],c_t[657],c_t2[658],s_t2[658]);
fa fau_1_659(b_i_s[659],s_t[659],c_t[658],c_t2[659],s_t2[659]);
fa fau_1_660(b_i_s[660],s_t[660],c_t[659],c_t2[660],s_t2[660]);
fa fau_1_661(b_i_s[661],s_t[661],c_t[660],c_t2[661],s_t2[661]);
fa fau_1_662(b_i_s[662],s_t[662],c_t[661],c_t2[662],s_t2[662]);
fa fau_1_663(b_i_s[663],s_t[663],c_t[662],c_t2[663],s_t2[663]);
fa fau_1_664(b_i_s[664],s_t[664],c_t[663],c_t2[664],s_t2[664]);
fa fau_1_665(b_i_s[665],s_t[665],c_t[664],c_t2[665],s_t2[665]);
fa fau_1_666(b_i_s[666],s_t[666],c_t[665],c_t2[666],s_t2[666]);
fa fau_1_667(b_i_s[667],s_t[667],c_t[666],c_t2[667],s_t2[667]);
fa fau_1_668(b_i_s[668],s_t[668],c_t[667],c_t2[668],s_t2[668]);
fa fau_1_669(b_i_s[669],s_t[669],c_t[668],c_t2[669],s_t2[669]);
fa fau_1_670(b_i_s[670],s_t[670],c_t[669],c_t2[670],s_t2[670]);
fa fau_1_671(b_i_s[671],s_t[671],c_t[670],c_t2[671],s_t2[671]);
fa fau_1_672(b_i_s[672],s_t[672],c_t[671],c_t2[672],s_t2[672]);
fa fau_1_673(b_i_s[673],s_t[673],c_t[672],c_t2[673],s_t2[673]);
fa fau_1_674(b_i_s[674],s_t[674],c_t[673],c_t2[674],s_t2[674]);
fa fau_1_675(b_i_s[675],s_t[675],c_t[674],c_t2[675],s_t2[675]);
fa fau_1_676(b_i_s[676],s_t[676],c_t[675],c_t2[676],s_t2[676]);
fa fau_1_677(b_i_s[677],s_t[677],c_t[676],c_t2[677],s_t2[677]);
fa fau_1_678(b_i_s[678],s_t[678],c_t[677],c_t2[678],s_t2[678]);
fa fau_1_679(b_i_s[679],s_t[679],c_t[678],c_t2[679],s_t2[679]);
fa fau_1_680(b_i_s[680],s_t[680],c_t[679],c_t2[680],s_t2[680]);
fa fau_1_681(b_i_s[681],s_t[681],c_t[680],c_t2[681],s_t2[681]);
fa fau_1_682(b_i_s[682],s_t[682],c_t[681],c_t2[682],s_t2[682]);
fa fau_1_683(b_i_s[683],s_t[683],c_t[682],c_t2[683],s_t2[683]);
fa fau_1_684(b_i_s[684],s_t[684],c_t[683],c_t2[684],s_t2[684]);
fa fau_1_685(b_i_s[685],s_t[685],c_t[684],c_t2[685],s_t2[685]);
fa fau_1_686(b_i_s[686],s_t[686],c_t[685],c_t2[686],s_t2[686]);
fa fau_1_687(b_i_s[687],s_t[687],c_t[686],c_t2[687],s_t2[687]);
fa fau_1_688(b_i_s[688],s_t[688],c_t[687],c_t2[688],s_t2[688]);
fa fau_1_689(b_i_s[689],s_t[689],c_t[688],c_t2[689],s_t2[689]);
fa fau_1_690(b_i_s[690],s_t[690],c_t[689],c_t2[690],s_t2[690]);
fa fau_1_691(b_i_s[691],s_t[691],c_t[690],c_t2[691],s_t2[691]);
fa fau_1_692(b_i_s[692],s_t[692],c_t[691],c_t2[692],s_t2[692]);
fa fau_1_693(b_i_s[693],s_t[693],c_t[692],c_t2[693],s_t2[693]);
fa fau_1_694(b_i_s[694],s_t[694],c_t[693],c_t2[694],s_t2[694]);
fa fau_1_695(b_i_s[695],s_t[695],c_t[694],c_t2[695],s_t2[695]);
fa fau_1_696(b_i_s[696],s_t[696],c_t[695],c_t2[696],s_t2[696]);
fa fau_1_697(b_i_s[697],s_t[697],c_t[696],c_t2[697],s_t2[697]);
fa fau_1_698(b_i_s[698],s_t[698],c_t[697],c_t2[698],s_t2[698]);
fa fau_1_699(b_i_s[699],s_t[699],c_t[698],c_t2[699],s_t2[699]);
fa fau_1_700(b_i_s[700],s_t[700],c_t[699],c_t2[700],s_t2[700]);
fa fau_1_701(b_i_s[701],s_t[701],c_t[700],c_t2[701],s_t2[701]);
fa fau_1_702(b_i_s[702],s_t[702],c_t[701],c_t2[702],s_t2[702]);
fa fau_1_703(b_i_s[703],s_t[703],c_t[702],c_t2[703],s_t2[703]);
fa fau_1_704(b_i_s[704],s_t[704],c_t[703],c_t2[704],s_t2[704]);
fa fau_1_705(b_i_s[705],s_t[705],c_t[704],c_t2[705],s_t2[705]);
fa fau_1_706(b_i_s[706],s_t[706],c_t[705],c_t2[706],s_t2[706]);
fa fau_1_707(b_i_s[707],s_t[707],c_t[706],c_t2[707],s_t2[707]);
fa fau_1_708(b_i_s[708],s_t[708],c_t[707],c_t2[708],s_t2[708]);
fa fau_1_709(b_i_s[709],s_t[709],c_t[708],c_t2[709],s_t2[709]);
fa fau_1_710(b_i_s[710],s_t[710],c_t[709],c_t2[710],s_t2[710]);
fa fau_1_711(b_i_s[711],s_t[711],c_t[710],c_t2[711],s_t2[711]);
fa fau_1_712(b_i_s[712],s_t[712],c_t[711],c_t2[712],s_t2[712]);
fa fau_1_713(b_i_s[713],s_t[713],c_t[712],c_t2[713],s_t2[713]);
fa fau_1_714(b_i_s[714],s_t[714],c_t[713],c_t2[714],s_t2[714]);
fa fau_1_715(b_i_s[715],s_t[715],c_t[714],c_t2[715],s_t2[715]);
fa fau_1_716(b_i_s[716],s_t[716],c_t[715],c_t2[716],s_t2[716]);
fa fau_1_717(b_i_s[717],s_t[717],c_t[716],c_t2[717],s_t2[717]);
fa fau_1_718(b_i_s[718],s_t[718],c_t[717],c_t2[718],s_t2[718]);
fa fau_1_719(b_i_s[719],s_t[719],c_t[718],c_t2[719],s_t2[719]);
fa fau_1_720(b_i_s[720],s_t[720],c_t[719],c_t2[720],s_t2[720]);
fa fau_1_721(b_i_s[721],s_t[721],c_t[720],c_t2[721],s_t2[721]);
fa fau_1_722(b_i_s[722],s_t[722],c_t[721],c_t2[722],s_t2[722]);
fa fau_1_723(b_i_s[723],s_t[723],c_t[722],c_t2[723],s_t2[723]);
fa fau_1_724(b_i_s[724],s_t[724],c_t[723],c_t2[724],s_t2[724]);
fa fau_1_725(b_i_s[725],s_t[725],c_t[724],c_t2[725],s_t2[725]);
fa fau_1_726(b_i_s[726],s_t[726],c_t[725],c_t2[726],s_t2[726]);
fa fau_1_727(b_i_s[727],s_t[727],c_t[726],c_t2[727],s_t2[727]);
fa fau_1_728(b_i_s[728],s_t[728],c_t[727],c_t2[728],s_t2[728]);
fa fau_1_729(b_i_s[729],s_t[729],c_t[728],c_t2[729],s_t2[729]);
fa fau_1_730(b_i_s[730],s_t[730],c_t[729],c_t2[730],s_t2[730]);
fa fau_1_731(b_i_s[731],s_t[731],c_t[730],c_t2[731],s_t2[731]);
fa fau_1_732(b_i_s[732],s_t[732],c_t[731],c_t2[732],s_t2[732]);
fa fau_1_733(b_i_s[733],s_t[733],c_t[732],c_t2[733],s_t2[733]);
fa fau_1_734(b_i_s[734],s_t[734],c_t[733],c_t2[734],s_t2[734]);
fa fau_1_735(b_i_s[735],s_t[735],c_t[734],c_t2[735],s_t2[735]);
fa fau_1_736(b_i_s[736],s_t[736],c_t[735],c_t2[736],s_t2[736]);
fa fau_1_737(b_i_s[737],s_t[737],c_t[736],c_t2[737],s_t2[737]);
fa fau_1_738(b_i_s[738],s_t[738],c_t[737],c_t2[738],s_t2[738]);
fa fau_1_739(b_i_s[739],s_t[739],c_t[738],c_t2[739],s_t2[739]);
fa fau_1_740(b_i_s[740],s_t[740],c_t[739],c_t2[740],s_t2[740]);
fa fau_1_741(b_i_s[741],s_t[741],c_t[740],c_t2[741],s_t2[741]);
fa fau_1_742(b_i_s[742],s_t[742],c_t[741],c_t2[742],s_t2[742]);
fa fau_1_743(b_i_s[743],s_t[743],c_t[742],c_t2[743],s_t2[743]);
fa fau_1_744(b_i_s[744],s_t[744],c_t[743],c_t2[744],s_t2[744]);
fa fau_1_745(b_i_s[745],s_t[745],c_t[744],c_t2[745],s_t2[745]);
fa fau_1_746(b_i_s[746],s_t[746],c_t[745],c_t2[746],s_t2[746]);
fa fau_1_747(b_i_s[747],s_t[747],c_t[746],c_t2[747],s_t2[747]);
fa fau_1_748(b_i_s[748],s_t[748],c_t[747],c_t2[748],s_t2[748]);
fa fau_1_749(b_i_s[749],s_t[749],c_t[748],c_t2[749],s_t2[749]);
fa fau_1_750(b_i_s[750],s_t[750],c_t[749],c_t2[750],s_t2[750]);
fa fau_1_751(b_i_s[751],s_t[751],c_t[750],c_t2[751],s_t2[751]);
fa fau_1_752(b_i_s[752],s_t[752],c_t[751],c_t2[752],s_t2[752]);
fa fau_1_753(b_i_s[753],s_t[753],c_t[752],c_t2[753],s_t2[753]);
fa fau_1_754(b_i_s[754],s_t[754],c_t[753],c_t2[754],s_t2[754]);
fa fau_1_755(b_i_s[755],s_t[755],c_t[754],c_t2[755],s_t2[755]);
fa fau_1_756(b_i_s[756],s_t[756],c_t[755],c_t2[756],s_t2[756]);
fa fau_1_757(b_i_s[757],s_t[757],c_t[756],c_t2[757],s_t2[757]);
fa fau_1_758(b_i_s[758],s_t[758],c_t[757],c_t2[758],s_t2[758]);
fa fau_1_759(b_i_s[759],s_t[759],c_t[758],c_t2[759],s_t2[759]);
fa fau_1_760(b_i_s[760],s_t[760],c_t[759],c_t2[760],s_t2[760]);
fa fau_1_761(b_i_s[761],s_t[761],c_t[760],c_t2[761],s_t2[761]);
fa fau_1_762(b_i_s[762],s_t[762],c_t[761],c_t2[762],s_t2[762]);
fa fau_1_763(b_i_s[763],s_t[763],c_t[762],c_t2[763],s_t2[763]);
fa fau_1_764(b_i_s[764],s_t[764],c_t[763],c_t2[764],s_t2[764]);
fa fau_1_765(b_i_s[765],s_t[765],c_t[764],c_t2[765],s_t2[765]);
fa fau_1_766(b_i_s[766],s_t[766],c_t[765],c_t2[766],s_t2[766]);
fa fau_1_767(b_i_s[767],s_t[767],c_t[766],c_t2[767],s_t2[767]);
fa fau_1_768(b_i_s[768],s_t[768],c_t[767],c_t2[768],s_t2[768]);
fa fau_1_769(b_i_s[769],s_t[769],c_t[768],c_t2[769],s_t2[769]);
fa fau_1_770(b_i_s[770],s_t[770],c_t[769],c_t2[770],s_t2[770]);
fa fau_1_771(b_i_s[771],s_t[771],c_t[770],c_t2[771],s_t2[771]);
fa fau_1_772(b_i_s[772],s_t[772],c_t[771],c_t2[772],s_t2[772]);
fa fau_1_773(b_i_s[773],s_t[773],c_t[772],c_t2[773],s_t2[773]);
fa fau_1_774(b_i_s[774],s_t[774],c_t[773],c_t2[774],s_t2[774]);
fa fau_1_775(b_i_s[775],s_t[775],c_t[774],c_t2[775],s_t2[775]);
fa fau_1_776(b_i_s[776],s_t[776],c_t[775],c_t2[776],s_t2[776]);
fa fau_1_777(b_i_s[777],s_t[777],c_t[776],c_t2[777],s_t2[777]);
fa fau_1_778(b_i_s[778],s_t[778],c_t[777],c_t2[778],s_t2[778]);
fa fau_1_779(b_i_s[779],s_t[779],c_t[778],c_t2[779],s_t2[779]);
fa fau_1_780(b_i_s[780],s_t[780],c_t[779],c_t2[780],s_t2[780]);
fa fau_1_781(b_i_s[781],s_t[781],c_t[780],c_t2[781],s_t2[781]);
fa fau_1_782(b_i_s[782],s_t[782],c_t[781],c_t2[782],s_t2[782]);
fa fau_1_783(b_i_s[783],s_t[783],c_t[782],c_t2[783],s_t2[783]);
fa fau_1_784(b_i_s[784],s_t[784],c_t[783],c_t2[784],s_t2[784]);
fa fau_1_785(b_i_s[785],s_t[785],c_t[784],c_t2[785],s_t2[785]);
fa fau_1_786(b_i_s[786],s_t[786],c_t[785],c_t2[786],s_t2[786]);
fa fau_1_787(b_i_s[787],s_t[787],c_t[786],c_t2[787],s_t2[787]);
fa fau_1_788(b_i_s[788],s_t[788],c_t[787],c_t2[788],s_t2[788]);
fa fau_1_789(b_i_s[789],s_t[789],c_t[788],c_t2[789],s_t2[789]);
fa fau_1_790(b_i_s[790],s_t[790],c_t[789],c_t2[790],s_t2[790]);
fa fau_1_791(b_i_s[791],s_t[791],c_t[790],c_t2[791],s_t2[791]);
fa fau_1_792(b_i_s[792],s_t[792],c_t[791],c_t2[792],s_t2[792]);
fa fau_1_793(b_i_s[793],s_t[793],c_t[792],c_t2[793],s_t2[793]);
fa fau_1_794(b_i_s[794],s_t[794],c_t[793],c_t2[794],s_t2[794]);
fa fau_1_795(b_i_s[795],s_t[795],c_t[794],c_t2[795],s_t2[795]);
fa fau_1_796(b_i_s[796],s_t[796],c_t[795],c_t2[796],s_t2[796]);
fa fau_1_797(b_i_s[797],s_t[797],c_t[796],c_t2[797],s_t2[797]);
fa fau_1_798(b_i_s[798],s_t[798],c_t[797],c_t2[798],s_t2[798]);
fa fau_1_799(b_i_s[799],s_t[799],c_t[798],c_t2[799],s_t2[799]);
fa fau_1_800(b_i_s[800],s_t[800],c_t[799],c_t2[800],s_t2[800]);
fa fau_1_801(b_i_s[801],s_t[801],c_t[800],c_t2[801],s_t2[801]);
fa fau_1_802(b_i_s[802],s_t[802],c_t[801],c_t2[802],s_t2[802]);
fa fau_1_803(b_i_s[803],s_t[803],c_t[802],c_t2[803],s_t2[803]);
fa fau_1_804(b_i_s[804],s_t[804],c_t[803],c_t2[804],s_t2[804]);
fa fau_1_805(b_i_s[805],s_t[805],c_t[804],c_t2[805],s_t2[805]);
fa fau_1_806(b_i_s[806],s_t[806],c_t[805],c_t2[806],s_t2[806]);
fa fau_1_807(b_i_s[807],s_t[807],c_t[806],c_t2[807],s_t2[807]);
fa fau_1_808(b_i_s[808],s_t[808],c_t[807],c_t2[808],s_t2[808]);
fa fau_1_809(b_i_s[809],s_t[809],c_t[808],c_t2[809],s_t2[809]);
fa fau_1_810(b_i_s[810],s_t[810],c_t[809],c_t2[810],s_t2[810]);
fa fau_1_811(b_i_s[811],s_t[811],c_t[810],c_t2[811],s_t2[811]);
fa fau_1_812(b_i_s[812],s_t[812],c_t[811],c_t2[812],s_t2[812]);
fa fau_1_813(b_i_s[813],s_t[813],c_t[812],c_t2[813],s_t2[813]);
fa fau_1_814(b_i_s[814],s_t[814],c_t[813],c_t2[814],s_t2[814]);
fa fau_1_815(b_i_s[815],s_t[815],c_t[814],c_t2[815],s_t2[815]);
fa fau_1_816(b_i_s[816],s_t[816],c_t[815],c_t2[816],s_t2[816]);
fa fau_1_817(b_i_s[817],s_t[817],c_t[816],c_t2[817],s_t2[817]);
fa fau_1_818(b_i_s[818],s_t[818],c_t[817],c_t2[818],s_t2[818]);
fa fau_1_819(b_i_s[819],s_t[819],c_t[818],c_t2[819],s_t2[819]);
fa fau_1_820(b_i_s[820],s_t[820],c_t[819],c_t2[820],s_t2[820]);
fa fau_1_821(b_i_s[821],s_t[821],c_t[820],c_t2[821],s_t2[821]);
fa fau_1_822(b_i_s[822],s_t[822],c_t[821],c_t2[822],s_t2[822]);
fa fau_1_823(b_i_s[823],s_t[823],c_t[822],c_t2[823],s_t2[823]);
fa fau_1_824(b_i_s[824],s_t[824],c_t[823],c_t2[824],s_t2[824]);
fa fau_1_825(b_i_s[825],s_t[825],c_t[824],c_t2[825],s_t2[825]);
fa fau_1_826(b_i_s[826],s_t[826],c_t[825],c_t2[826],s_t2[826]);
fa fau_1_827(b_i_s[827],s_t[827],c_t[826],c_t2[827],s_t2[827]);
fa fau_1_828(b_i_s[828],s_t[828],c_t[827],c_t2[828],s_t2[828]);
fa fau_1_829(b_i_s[829],s_t[829],c_t[828],c_t2[829],s_t2[829]);
fa fau_1_830(b_i_s[830],s_t[830],c_t[829],c_t2[830],s_t2[830]);
fa fau_1_831(b_i_s[831],s_t[831],c_t[830],c_t2[831],s_t2[831]);
fa fau_1_832(b_i_s[832],s_t[832],c_t[831],c_t2[832],s_t2[832]);
fa fau_1_833(b_i_s[833],s_t[833],c_t[832],c_t2[833],s_t2[833]);
fa fau_1_834(b_i_s[834],s_t[834],c_t[833],c_t2[834],s_t2[834]);
fa fau_1_835(b_i_s[835],s_t[835],c_t[834],c_t2[835],s_t2[835]);
fa fau_1_836(b_i_s[836],s_t[836],c_t[835],c_t2[836],s_t2[836]);
fa fau_1_837(b_i_s[837],s_t[837],c_t[836],c_t2[837],s_t2[837]);
fa fau_1_838(b_i_s[838],s_t[838],c_t[837],c_t2[838],s_t2[838]);
fa fau_1_839(b_i_s[839],s_t[839],c_t[838],c_t2[839],s_t2[839]);
fa fau_1_840(b_i_s[840],s_t[840],c_t[839],c_t2[840],s_t2[840]);
fa fau_1_841(b_i_s[841],s_t[841],c_t[840],c_t2[841],s_t2[841]);
fa fau_1_842(b_i_s[842],s_t[842],c_t[841],c_t2[842],s_t2[842]);
fa fau_1_843(b_i_s[843],s_t[843],c_t[842],c_t2[843],s_t2[843]);
fa fau_1_844(b_i_s[844],s_t[844],c_t[843],c_t2[844],s_t2[844]);
fa fau_1_845(b_i_s[845],s_t[845],c_t[844],c_t2[845],s_t2[845]);
fa fau_1_846(b_i_s[846],s_t[846],c_t[845],c_t2[846],s_t2[846]);
fa fau_1_847(b_i_s[847],s_t[847],c_t[846],c_t2[847],s_t2[847]);
fa fau_1_848(b_i_s[848],s_t[848],c_t[847],c_t2[848],s_t2[848]);
fa fau_1_849(b_i_s[849],s_t[849],c_t[848],c_t2[849],s_t2[849]);
fa fau_1_850(b_i_s[850],s_t[850],c_t[849],c_t2[850],s_t2[850]);
fa fau_1_851(b_i_s[851],s_t[851],c_t[850],c_t2[851],s_t2[851]);
fa fau_1_852(b_i_s[852],s_t[852],c_t[851],c_t2[852],s_t2[852]);
fa fau_1_853(b_i_s[853],s_t[853],c_t[852],c_t2[853],s_t2[853]);
fa fau_1_854(b_i_s[854],s_t[854],c_t[853],c_t2[854],s_t2[854]);
fa fau_1_855(b_i_s[855],s_t[855],c_t[854],c_t2[855],s_t2[855]);
fa fau_1_856(b_i_s[856],s_t[856],c_t[855],c_t2[856],s_t2[856]);
fa fau_1_857(b_i_s[857],s_t[857],c_t[856],c_t2[857],s_t2[857]);
fa fau_1_858(b_i_s[858],s_t[858],c_t[857],c_t2[858],s_t2[858]);
fa fau_1_859(b_i_s[859],s_t[859],c_t[858],c_t2[859],s_t2[859]);
fa fau_1_860(b_i_s[860],s_t[860],c_t[859],c_t2[860],s_t2[860]);
fa fau_1_861(b_i_s[861],s_t[861],c_t[860],c_t2[861],s_t2[861]);
fa fau_1_862(b_i_s[862],s_t[862],c_t[861],c_t2[862],s_t2[862]);
fa fau_1_863(b_i_s[863],s_t[863],c_t[862],c_t2[863],s_t2[863]);
fa fau_1_864(b_i_s[864],s_t[864],c_t[863],c_t2[864],s_t2[864]);
fa fau_1_865(b_i_s[865],s_t[865],c_t[864],c_t2[865],s_t2[865]);
fa fau_1_866(b_i_s[866],s_t[866],c_t[865],c_t2[866],s_t2[866]);
fa fau_1_867(b_i_s[867],s_t[867],c_t[866],c_t2[867],s_t2[867]);
fa fau_1_868(b_i_s[868],s_t[868],c_t[867],c_t2[868],s_t2[868]);
fa fau_1_869(b_i_s[869],s_t[869],c_t[868],c_t2[869],s_t2[869]);
fa fau_1_870(b_i_s[870],s_t[870],c_t[869],c_t2[870],s_t2[870]);
fa fau_1_871(b_i_s[871],s_t[871],c_t[870],c_t2[871],s_t2[871]);
fa fau_1_872(b_i_s[872],s_t[872],c_t[871],c_t2[872],s_t2[872]);
fa fau_1_873(b_i_s[873],s_t[873],c_t[872],c_t2[873],s_t2[873]);
fa fau_1_874(b_i_s[874],s_t[874],c_t[873],c_t2[874],s_t2[874]);
fa fau_1_875(b_i_s[875],s_t[875],c_t[874],c_t2[875],s_t2[875]);
fa fau_1_876(b_i_s[876],s_t[876],c_t[875],c_t2[876],s_t2[876]);
fa fau_1_877(b_i_s[877],s_t[877],c_t[876],c_t2[877],s_t2[877]);
fa fau_1_878(b_i_s[878],s_t[878],c_t[877],c_t2[878],s_t2[878]);
fa fau_1_879(b_i_s[879],s_t[879],c_t[878],c_t2[879],s_t2[879]);
fa fau_1_880(b_i_s[880],s_t[880],c_t[879],c_t2[880],s_t2[880]);
fa fau_1_881(b_i_s[881],s_t[881],c_t[880],c_t2[881],s_t2[881]);
fa fau_1_882(b_i_s[882],s_t[882],c_t[881],c_t2[882],s_t2[882]);
fa fau_1_883(b_i_s[883],s_t[883],c_t[882],c_t2[883],s_t2[883]);
fa fau_1_884(b_i_s[884],s_t[884],c_t[883],c_t2[884],s_t2[884]);
fa fau_1_885(b_i_s[885],s_t[885],c_t[884],c_t2[885],s_t2[885]);
fa fau_1_886(b_i_s[886],s_t[886],c_t[885],c_t2[886],s_t2[886]);
fa fau_1_887(b_i_s[887],s_t[887],c_t[886],c_t2[887],s_t2[887]);
fa fau_1_888(b_i_s[888],s_t[888],c_t[887],c_t2[888],s_t2[888]);
fa fau_1_889(b_i_s[889],s_t[889],c_t[888],c_t2[889],s_t2[889]);
fa fau_1_890(b_i_s[890],s_t[890],c_t[889],c_t2[890],s_t2[890]);
fa fau_1_891(b_i_s[891],s_t[891],c_t[890],c_t2[891],s_t2[891]);
fa fau_1_892(b_i_s[892],s_t[892],c_t[891],c_t2[892],s_t2[892]);
fa fau_1_893(b_i_s[893],s_t[893],c_t[892],c_t2[893],s_t2[893]);
fa fau_1_894(b_i_s[894],s_t[894],c_t[893],c_t2[894],s_t2[894]);
fa fau_1_895(b_i_s[895],s_t[895],c_t[894],c_t2[895],s_t2[895]);
fa fau_1_896(b_i_s[896],s_t[896],c_t[895],c_t2[896],s_t2[896]);
fa fau_1_897(b_i_s[897],s_t[897],c_t[896],c_t2[897],s_t2[897]);
fa fau_1_898(b_i_s[898],s_t[898],c_t[897],c_t2[898],s_t2[898]);
fa fau_1_899(b_i_s[899],s_t[899],c_t[898],c_t2[899],s_t2[899]);
fa fau_1_900(b_i_s[900],s_t[900],c_t[899],c_t2[900],s_t2[900]);
fa fau_1_901(b_i_s[901],s_t[901],c_t[900],c_t2[901],s_t2[901]);
fa fau_1_902(b_i_s[902],s_t[902],c_t[901],c_t2[902],s_t2[902]);
fa fau_1_903(b_i_s[903],s_t[903],c_t[902],c_t2[903],s_t2[903]);
fa fau_1_904(b_i_s[904],s_t[904],c_t[903],c_t2[904],s_t2[904]);
fa fau_1_905(b_i_s[905],s_t[905],c_t[904],c_t2[905],s_t2[905]);
fa fau_1_906(b_i_s[906],s_t[906],c_t[905],c_t2[906],s_t2[906]);
fa fau_1_907(b_i_s[907],s_t[907],c_t[906],c_t2[907],s_t2[907]);
fa fau_1_908(b_i_s[908],s_t[908],c_t[907],c_t2[908],s_t2[908]);
fa fau_1_909(b_i_s[909],s_t[909],c_t[908],c_t2[909],s_t2[909]);
fa fau_1_910(b_i_s[910],s_t[910],c_t[909],c_t2[910],s_t2[910]);
fa fau_1_911(b_i_s[911],s_t[911],c_t[910],c_t2[911],s_t2[911]);
fa fau_1_912(b_i_s[912],s_t[912],c_t[911],c_t2[912],s_t2[912]);
fa fau_1_913(b_i_s[913],s_t[913],c_t[912],c_t2[913],s_t2[913]);
fa fau_1_914(b_i_s[914],s_t[914],c_t[913],c_t2[914],s_t2[914]);
fa fau_1_915(b_i_s[915],s_t[915],c_t[914],c_t2[915],s_t2[915]);
fa fau_1_916(b_i_s[916],s_t[916],c_t[915],c_t2[916],s_t2[916]);
fa fau_1_917(b_i_s[917],s_t[917],c_t[916],c_t2[917],s_t2[917]);
fa fau_1_918(b_i_s[918],s_t[918],c_t[917],c_t2[918],s_t2[918]);
fa fau_1_919(b_i_s[919],s_t[919],c_t[918],c_t2[919],s_t2[919]);
fa fau_1_920(b_i_s[920],s_t[920],c_t[919],c_t2[920],s_t2[920]);
fa fau_1_921(b_i_s[921],s_t[921],c_t[920],c_t2[921],s_t2[921]);
fa fau_1_922(b_i_s[922],s_t[922],c_t[921],c_t2[922],s_t2[922]);
fa fau_1_923(b_i_s[923],s_t[923],c_t[922],c_t2[923],s_t2[923]);
fa fau_1_924(b_i_s[924],s_t[924],c_t[923],c_t2[924],s_t2[924]);
fa fau_1_925(b_i_s[925],s_t[925],c_t[924],c_t2[925],s_t2[925]);
fa fau_1_926(b_i_s[926],s_t[926],c_t[925],c_t2[926],s_t2[926]);
fa fau_1_927(b_i_s[927],s_t[927],c_t[926],c_t2[927],s_t2[927]);
fa fau_1_928(b_i_s[928],s_t[928],c_t[927],c_t2[928],s_t2[928]);
fa fau_1_929(b_i_s[929],s_t[929],c_t[928],c_t2[929],s_t2[929]);
fa fau_1_930(b_i_s[930],s_t[930],c_t[929],c_t2[930],s_t2[930]);
fa fau_1_931(b_i_s[931],s_t[931],c_t[930],c_t2[931],s_t2[931]);
fa fau_1_932(b_i_s[932],s_t[932],c_t[931],c_t2[932],s_t2[932]);
fa fau_1_933(b_i_s[933],s_t[933],c_t[932],c_t2[933],s_t2[933]);
fa fau_1_934(b_i_s[934],s_t[934],c_t[933],c_t2[934],s_t2[934]);
fa fau_1_935(b_i_s[935],s_t[935],c_t[934],c_t2[935],s_t2[935]);
fa fau_1_936(b_i_s[936],s_t[936],c_t[935],c_t2[936],s_t2[936]);
fa fau_1_937(b_i_s[937],s_t[937],c_t[936],c_t2[937],s_t2[937]);
fa fau_1_938(b_i_s[938],s_t[938],c_t[937],c_t2[938],s_t2[938]);
fa fau_1_939(b_i_s[939],s_t[939],c_t[938],c_t2[939],s_t2[939]);
fa fau_1_940(b_i_s[940],s_t[940],c_t[939],c_t2[940],s_t2[940]);
fa fau_1_941(b_i_s[941],s_t[941],c_t[940],c_t2[941],s_t2[941]);
fa fau_1_942(b_i_s[942],s_t[942],c_t[941],c_t2[942],s_t2[942]);
fa fau_1_943(b_i_s[943],s_t[943],c_t[942],c_t2[943],s_t2[943]);
fa fau_1_944(b_i_s[944],s_t[944],c_t[943],c_t2[944],s_t2[944]);
fa fau_1_945(b_i_s[945],s_t[945],c_t[944],c_t2[945],s_t2[945]);
fa fau_1_946(b_i_s[946],s_t[946],c_t[945],c_t2[946],s_t2[946]);
fa fau_1_947(b_i_s[947],s_t[947],c_t[946],c_t2[947],s_t2[947]);
fa fau_1_948(b_i_s[948],s_t[948],c_t[947],c_t2[948],s_t2[948]);
fa fau_1_949(b_i_s[949],s_t[949],c_t[948],c_t2[949],s_t2[949]);
fa fau_1_950(b_i_s[950],s_t[950],c_t[949],c_t2[950],s_t2[950]);
fa fau_1_951(b_i_s[951],s_t[951],c_t[950],c_t2[951],s_t2[951]);
fa fau_1_952(b_i_s[952],s_t[952],c_t[951],c_t2[952],s_t2[952]);
fa fau_1_953(b_i_s[953],s_t[953],c_t[952],c_t2[953],s_t2[953]);
fa fau_1_954(b_i_s[954],s_t[954],c_t[953],c_t2[954],s_t2[954]);
fa fau_1_955(b_i_s[955],s_t[955],c_t[954],c_t2[955],s_t2[955]);
fa fau_1_956(b_i_s[956],s_t[956],c_t[955],c_t2[956],s_t2[956]);
fa fau_1_957(b_i_s[957],s_t[957],c_t[956],c_t2[957],s_t2[957]);
fa fau_1_958(b_i_s[958],s_t[958],c_t[957],c_t2[958],s_t2[958]);
fa fau_1_959(b_i_s[959],s_t[959],c_t[958],c_t2[959],s_t2[959]);
fa fau_1_960(b_i_s[960],s_t[960],c_t[959],c_t2[960],s_t2[960]);
fa fau_1_961(b_i_s[961],s_t[961],c_t[960],c_t2[961],s_t2[961]);
fa fau_1_962(b_i_s[962],s_t[962],c_t[961],c_t2[962],s_t2[962]);
fa fau_1_963(b_i_s[963],s_t[963],c_t[962],c_t2[963],s_t2[963]);
fa fau_1_964(b_i_s[964],s_t[964],c_t[963],c_t2[964],s_t2[964]);
fa fau_1_965(b_i_s[965],s_t[965],c_t[964],c_t2[965],s_t2[965]);
fa fau_1_966(b_i_s[966],s_t[966],c_t[965],c_t2[966],s_t2[966]);
fa fau_1_967(b_i_s[967],s_t[967],c_t[966],c_t2[967],s_t2[967]);
fa fau_1_968(b_i_s[968],s_t[968],c_t[967],c_t2[968],s_t2[968]);
fa fau_1_969(b_i_s[969],s_t[969],c_t[968],c_t2[969],s_t2[969]);
fa fau_1_970(b_i_s[970],s_t[970],c_t[969],c_t2[970],s_t2[970]);
fa fau_1_971(b_i_s[971],s_t[971],c_t[970],c_t2[971],s_t2[971]);
fa fau_1_972(b_i_s[972],s_t[972],c_t[971],c_t2[972],s_t2[972]);
fa fau_1_973(b_i_s[973],s_t[973],c_t[972],c_t2[973],s_t2[973]);
fa fau_1_974(b_i_s[974],s_t[974],c_t[973],c_t2[974],s_t2[974]);
fa fau_1_975(b_i_s[975],s_t[975],c_t[974],c_t2[975],s_t2[975]);
fa fau_1_976(b_i_s[976],s_t[976],c_t[975],c_t2[976],s_t2[976]);
fa fau_1_977(b_i_s[977],s_t[977],c_t[976],c_t2[977],s_t2[977]);
fa fau_1_978(b_i_s[978],s_t[978],c_t[977],c_t2[978],s_t2[978]);
fa fau_1_979(b_i_s[979],s_t[979],c_t[978],c_t2[979],s_t2[979]);
fa fau_1_980(b_i_s[980],s_t[980],c_t[979],c_t2[980],s_t2[980]);
fa fau_1_981(b_i_s[981],s_t[981],c_t[980],c_t2[981],s_t2[981]);
fa fau_1_982(b_i_s[982],s_t[982],c_t[981],c_t2[982],s_t2[982]);
fa fau_1_983(b_i_s[983],s_t[983],c_t[982],c_t2[983],s_t2[983]);
fa fau_1_984(b_i_s[984],s_t[984],c_t[983],c_t2[984],s_t2[984]);
fa fau_1_985(b_i_s[985],s_t[985],c_t[984],c_t2[985],s_t2[985]);
fa fau_1_986(b_i_s[986],s_t[986],c_t[985],c_t2[986],s_t2[986]);
fa fau_1_987(b_i_s[987],s_t[987],c_t[986],c_t2[987],s_t2[987]);
fa fau_1_988(b_i_s[988],s_t[988],c_t[987],c_t2[988],s_t2[988]);
fa fau_1_989(b_i_s[989],s_t[989],c_t[988],c_t2[989],s_t2[989]);
fa fau_1_990(b_i_s[990],s_t[990],c_t[989],c_t2[990],s_t2[990]);
fa fau_1_991(b_i_s[991],s_t[991],c_t[990],c_t2[991],s_t2[991]);
fa fau_1_992(b_i_s[992],s_t[992],c_t[991],c_t2[992],s_t2[992]);
fa fau_1_993(b_i_s[993],s_t[993],c_t[992],c_t2[993],s_t2[993]);
fa fau_1_994(b_i_s[994],s_t[994],c_t[993],c_t2[994],s_t2[994]);
fa fau_1_995(b_i_s[995],s_t[995],c_t[994],c_t2[995],s_t2[995]);
fa fau_1_996(b_i_s[996],s_t[996],c_t[995],c_t2[996],s_t2[996]);
fa fau_1_997(b_i_s[997],s_t[997],c_t[996],c_t2[997],s_t2[997]);
fa fau_1_998(b_i_s[998],s_t[998],c_t[997],c_t2[998],s_t2[998]);
fa fau_1_999(b_i_s[999],s_t[999],c_t[998],c_t2[999],s_t2[999]);
fa fau_1_1000(b_i_s[1000],s_t[1000],c_t[999],c_t2[1000],s_t2[1000]);
fa fau_1_1001(b_i_s[1001],s_t[1001],c_t[1000],c_t2[1001],s_t2[1001]);
fa fau_1_1002(b_i_s[1002],s_t[1002],c_t[1001],c_t2[1002],s_t2[1002]);
fa fau_1_1003(b_i_s[1003],s_t[1003],c_t[1002],c_t2[1003],s_t2[1003]);
fa fau_1_1004(b_i_s[1004],s_t[1004],c_t[1003],c_t2[1004],s_t2[1004]);
fa fau_1_1005(b_i_s[1005],s_t[1005],c_t[1004],c_t2[1005],s_t2[1005]);
fa fau_1_1006(b_i_s[1006],s_t[1006],c_t[1005],c_t2[1006],s_t2[1006]);
fa fau_1_1007(b_i_s[1007],s_t[1007],c_t[1006],c_t2[1007],s_t2[1007]);
fa fau_1_1008(b_i_s[1008],s_t[1008],c_t[1007],c_t2[1008],s_t2[1008]);
fa fau_1_1009(b_i_s[1009],s_t[1009],c_t[1008],c_t2[1009],s_t2[1009]);
fa fau_1_1010(b_i_s[1010],s_t[1010],c_t[1009],c_t2[1010],s_t2[1010]);
fa fau_1_1011(b_i_s[1011],s_t[1011],c_t[1010],c_t2[1011],s_t2[1011]);
fa fau_1_1012(b_i_s[1012],s_t[1012],c_t[1011],c_t2[1012],s_t2[1012]);
fa fau_1_1013(b_i_s[1013],s_t[1013],c_t[1012],c_t2[1013],s_t2[1013]);
fa fau_1_1014(b_i_s[1014],s_t[1014],c_t[1013],c_t2[1014],s_t2[1014]);
fa fau_1_1015(b_i_s[1015],s_t[1015],c_t[1014],c_t2[1015],s_t2[1015]);
fa fau_1_1016(b_i_s[1016],s_t[1016],c_t[1015],c_t2[1016],s_t2[1016]);
fa fau_1_1017(b_i_s[1017],s_t[1017],c_t[1016],c_t2[1017],s_t2[1017]);
fa fau_1_1018(b_i_s[1018],s_t[1018],c_t[1017],c_t2[1018],s_t2[1018]);
fa fau_1_1019(b_i_s[1019],s_t[1019],c_t[1018],c_t2[1019],s_t2[1019]);
fa fau_1_1020(b_i_s[1020],s_t[1020],c_t[1019],c_t2[1020],s_t2[1020]);
fa fau_1_1021(b_i_s[1021],s_t[1021],c_t[1020],c_t2[1021],s_t2[1021]);
fa fau_1_1022(b_i_s[1022],s_t[1022],c_t[1021],c_t2[1022],s_t2[1022]);
fa fau_1_1023(b_i_s[1023],s_t[1023],c_t[1022],c_t2[1023],s_t2[1023]);
fa fau_1_1024(b_i_s[1024],s_t[1024],c_t[1023],c_t2[1024],s_t2[1024]);
fa fau_1_1025(b_i_s[1025],s_t[1025],c_t[1024],c_t2[1025],s_t2[1025]);
fa fau_1_1026(b_i_s[1026],s_t[1026],c_t[1025],c_t2[1026],s_t2[1026]);
fa fau_1_1027(b_i_s[1027],s_t[1027],c_t[1026],c_t2[1027],s_t2[1027]);
fa fau_1_1028(b_i_s[1028],s_t[1028],c_t[1027],c_t2[1028],s_t2[1028]);
fa fau_1_1029(b_i_s[1029],s_t[1029],c_t[1028],c_t2[1029],s_t2[1029]);
fa fau_1_1030(b_i_s[1030],s_t[1030],c_t[1029],c_t2[1030],s_t2[1030]);
fa fau_1_1031(b_i_s[1031],s_t[1031],c_t[1030],c_t2[1031],s_t2[1031]);
fa fau_1_1032(b_i_s[1032],s_t[1032],c_t[1031],c_t2[1032],s_t2[1032]);
fa fau_1_1033(b_i_s[1033],s_t[1033],c_t[1032],c_t2[1033],s_t2[1033]);
fa fau_1_1034(b_i_s[1034],s_t[1034],c_t[1033],c_t2[1034],s_t2[1034]);
fa fau_1_1035(b_i_s[1035],s_t[1035],c_t[1034],c_t2[1035],s_t2[1035]);
fa fau_1_1036(b_i_s[1036],s_t[1036],c_t[1035],c_t2[1036],s_t2[1036]);
fa fau_1_1037(b_i_s[1037],s_t[1037],c_t[1036],c_t2[1037],s_t2[1037]);
fa fau_1_1038(b_i_s[1038],s_t[1038],c_t[1037],c_t2[1038],s_t2[1038]);
fa fau_1_1039(b_i_s[1039],s_t[1039],c_t[1038],c_t2[1039],s_t2[1039]);
fa fau_1_1040(b_i_s[1040],s_t[1040],c_t[1039],c_t2[1040],s_t2[1040]);
fa fau_1_1041(b_i_s[1041],s_t[1041],c_t[1040],c_t2[1041],s_t2[1041]);
fa fau_1_1042(b_i_s[1042],s_t[1042],c_t[1041],c_t2[1042],s_t2[1042]);
fa fau_1_1043(b_i_s[1043],s_t[1043],c_t[1042],c_t2[1043],s_t2[1043]);
fa fau_1_1044(b_i_s[1044],s_t[1044],c_t[1043],c_t2[1044],s_t2[1044]);
fa fau_1_1045(b_i_s[1045],s_t[1045],c_t[1044],c_t2[1045],s_t2[1045]);
fa fau_1_1046(b_i_s[1046],s_t[1046],c_t[1045],c_t2[1046],s_t2[1046]);
fa fau_1_1047(b_i_s[1047],s_t[1047],c_t[1046],c_t2[1047],s_t2[1047]);
fa fau_1_1048(b_i_s[1048],s_t[1048],c_t[1047],c_t2[1048],s_t2[1048]);
fa fau_1_1049(b_i_s[1049],s_t[1049],c_t[1048],c_t2[1049],s_t2[1049]);
fa fau_1_1050(b_i_s[1050],s_t[1050],c_t[1049],c_t2[1050],s_t2[1050]);
fa fau_1_1051(b_i_s[1051],s_t[1051],c_t[1050],c_t2[1051],s_t2[1051]);
fa fau_1_1052(b_i_s[1052],s_t[1052],c_t[1051],c_t2[1052],s_t2[1052]);
fa fau_1_1053(b_i_s[1053],s_t[1053],c_t[1052],c_t2[1053],s_t2[1053]);
fa fau_1_1054(b_i_s[1054],s_t[1054],c_t[1053],c_t2[1054],s_t2[1054]);
fa fau_1_1055(b_i_s[1055],s_t[1055],c_t[1054],c_t2[1055],s_t2[1055]);
fa fau_1_1056(b_i_s[1056],s_t[1056],c_t[1055],c_t2[1056],s_t2[1056]);
fa fau_1_1057(b_i_s[1057],s_t[1057],c_t[1056],c_t2[1057],s_t2[1057]);
fa fau_1_1058(b_i_s[1058],s_t[1058],c_t[1057],c_t2[1058],s_t2[1058]);
fa fau_1_1059(b_i_s[1059],s_t[1059],c_t[1058],c_t2[1059],s_t2[1059]);
fa fau_1_1060(b_i_s[1060],s_t[1060],c_t[1059],c_t2[1060],s_t2[1060]);
fa fau_1_1061(b_i_s[1061],s_t[1061],c_t[1060],c_t2[1061],s_t2[1061]);
fa fau_1_1062(b_i_s[1062],s_t[1062],c_t[1061],c_t2[1062],s_t2[1062]);
fa fau_1_1063(b_i_s[1063],s_t[1063],c_t[1062],c_t2[1063],s_t2[1063]);
fa fau_1_1064(b_i_s[1064],s_t[1064],c_t[1063],c_t2[1064],s_t2[1064]);
fa fau_1_1065(b_i_s[1065],s_t[1065],c_t[1064],c_t2[1065],s_t2[1065]);
fa fau_1_1066(b_i_s[1066],s_t[1066],c_t[1065],c_t2[1066],s_t2[1066]);
fa fau_1_1067(b_i_s[1067],s_t[1067],c_t[1066],c_t2[1067],s_t2[1067]);
fa fau_1_1068(b_i_s[1068],s_t[1068],c_t[1067],c_t2[1068],s_t2[1068]);
fa fau_1_1069(b_i_s[1069],s_t[1069],c_t[1068],c_t2[1069],s_t2[1069]);
fa fau_1_1070(b_i_s[1070],s_t[1070],c_t[1069],c_t2[1070],s_t2[1070]);
fa fau_1_1071(b_i_s[1071],s_t[1071],c_t[1070],c_t2[1071],s_t2[1071]);
fa fau_1_1072(b_i_s[1072],s_t[1072],c_t[1071],c_t2[1072],s_t2[1072]);
fa fau_1_1073(b_i_s[1073],s_t[1073],c_t[1072],c_t2[1073],s_t2[1073]);
fa fau_1_1074(b_i_s[1074],s_t[1074],c_t[1073],c_t2[1074],s_t2[1074]);
fa fau_1_1075(b_i_s[1075],s_t[1075],c_t[1074],c_t2[1075],s_t2[1075]);
fa fau_1_1076(b_i_s[1076],s_t[1076],c_t[1075],c_t2[1076],s_t2[1076]);
fa fau_1_1077(b_i_s[1077],s_t[1077],c_t[1076],c_t2[1077],s_t2[1077]);
fa fau_1_1078(b_i_s[1078],s_t[1078],c_t[1077],c_t2[1078],s_t2[1078]);
fa fau_1_1079(b_i_s[1079],s_t[1079],c_t[1078],c_t2[1079],s_t2[1079]);
fa fau_1_1080(b_i_s[1080],s_t[1080],c_t[1079],c_t2[1080],s_t2[1080]);
fa fau_1_1081(b_i_s[1081],s_t[1081],c_t[1080],c_t2[1081],s_t2[1081]);
fa fau_1_1082(b_i_s[1082],s_t[1082],c_t[1081],c_t2[1082],s_t2[1082]);
fa fau_1_1083(b_i_s[1083],s_t[1083],c_t[1082],c_t2[1083],s_t2[1083]);
fa fau_1_1084(b_i_s[1084],s_t[1084],c_t[1083],c_t2[1084],s_t2[1084]);
fa fau_1_1085(b_i_s[1085],s_t[1085],c_t[1084],c_t2[1085],s_t2[1085]);
fa fau_1_1086(b_i_s[1086],s_t[1086],c_t[1085],c_t2[1086],s_t2[1086]);
fa fau_1_1087(b_i_s[1087],s_t[1087],c_t[1086],c_t2[1087],s_t2[1087]);
fa fau_1_1088(b_i_s[1088],s_t[1088],c_t[1087],c_t2[1088],s_t2[1088]);
fa fau_1_1089(b_i_s[1089],s_t[1089],c_t[1088],c_t2[1089],s_t2[1089]);
fa fau_1_1090(b_i_s[1090],s_t[1090],c_t[1089],c_t2[1090],s_t2[1090]);
fa fau_1_1091(b_i_s[1091],s_t[1091],c_t[1090],c_t2[1091],s_t2[1091]);
fa fau_1_1092(b_i_s[1092],s_t[1092],c_t[1091],c_t2[1092],s_t2[1092]);
fa fau_1_1093(b_i_s[1093],s_t[1093],c_t[1092],c_t2[1093],s_t2[1093]);
fa fau_1_1094(b_i_s[1094],s_t[1094],c_t[1093],c_t2[1094],s_t2[1094]);
fa fau_1_1095(b_i_s[1095],s_t[1095],c_t[1094],c_t2[1095],s_t2[1095]);
fa fau_1_1096(b_i_s[1096],s_t[1096],c_t[1095],c_t2[1096],s_t2[1096]);
fa fau_1_1097(b_i_s[1097],s_t[1097],c_t[1096],c_t2[1097],s_t2[1097]);
fa fau_1_1098(b_i_s[1098],s_t[1098],c_t[1097],c_t2[1098],s_t2[1098]);
fa fau_1_1099(b_i_s[1099],s_t[1099],c_t[1098],c_t2[1099],s_t2[1099]);
fa fau_1_1100(b_i_s[1100],s_t[1100],c_t[1099],c_t2[1100],s_t2[1100]);
fa fau_1_1101(b_i_s[1101],s_t[1101],c_t[1100],c_t2[1101],s_t2[1101]);
fa fau_1_1102(b_i_s[1102],s_t[1102],c_t[1101],c_t2[1102],s_t2[1102]);
fa fau_1_1103(b_i_s[1103],s_t[1103],c_t[1102],c_t2[1103],s_t2[1103]);
fa fau_1_1104(b_i_s[1104],s_t[1104],c_t[1103],c_t2[1104],s_t2[1104]);
fa fau_1_1105(b_i_s[1105],s_t[1105],c_t[1104],c_t2[1105],s_t2[1105]);
fa fau_1_1106(b_i_s[1106],s_t[1106],c_t[1105],c_t2[1106],s_t2[1106]);
fa fau_1_1107(b_i_s[1107],s_t[1107],c_t[1106],c_t2[1107],s_t2[1107]);
fa fau_1_1108(b_i_s[1108],s_t[1108],c_t[1107],c_t2[1108],s_t2[1108]);
fa fau_1_1109(b_i_s[1109],s_t[1109],c_t[1108],c_t2[1109],s_t2[1109]);
fa fau_1_1110(b_i_s[1110],s_t[1110],c_t[1109],c_t2[1110],s_t2[1110]);
fa fau_1_1111(b_i_s[1111],s_t[1111],c_t[1110],c_t2[1111],s_t2[1111]);
fa fau_1_1112(b_i_s[1112],s_t[1112],c_t[1111],c_t2[1112],s_t2[1112]);
fa fau_1_1113(b_i_s[1113],s_t[1113],c_t[1112],c_t2[1113],s_t2[1113]);
fa fau_1_1114(b_i_s[1114],s_t[1114],c_t[1113],c_t2[1114],s_t2[1114]);
fa fau_1_1115(b_i_s[1115],s_t[1115],c_t[1114],c_t2[1115],s_t2[1115]);
fa fau_1_1116(b_i_s[1116],s_t[1116],c_t[1115],c_t2[1116],s_t2[1116]);
fa fau_1_1117(b_i_s[1117],s_t[1117],c_t[1116],c_t2[1117],s_t2[1117]);
fa fau_1_1118(b_i_s[1118],s_t[1118],c_t[1117],c_t2[1118],s_t2[1118]);
fa fau_1_1119(b_i_s[1119],s_t[1119],c_t[1118],c_t2[1119],s_t2[1119]);
fa fau_1_1120(b_i_s[1120],s_t[1120],c_t[1119],c_t2[1120],s_t2[1120]);
fa fau_1_1121(b_i_s[1121],s_t[1121],c_t[1120],c_t2[1121],s_t2[1121]);
fa fau_1_1122(b_i_s[1122],s_t[1122],c_t[1121],c_t2[1122],s_t2[1122]);
fa fau_1_1123(b_i_s[1123],s_t[1123],c_t[1122],c_t2[1123],s_t2[1123]);
fa fau_1_1124(b_i_s[1124],s_t[1124],c_t[1123],c_t2[1124],s_t2[1124]);
fa fau_1_1125(b_i_s[1125],s_t[1125],c_t[1124],c_t2[1125],s_t2[1125]);
fa fau_1_1126(b_i_s[1126],s_t[1126],c_t[1125],c_t2[1126],s_t2[1126]);
fa fau_1_1127(b_i_s[1127],s_t[1127],c_t[1126],c_t2[1127],s_t2[1127]);
fa fau_1_1128(b_i_s[1128],s_t[1128],c_t[1127],c_t2[1128],s_t2[1128]);
fa fau_1_1129(b_i_s[1129],s_t[1129],c_t[1128],c_t2[1129],s_t2[1129]);
fa fau_1_1130(b_i_s[1130],s_t[1130],c_t[1129],c_t2[1130],s_t2[1130]);
fa fau_1_1131(b_i_s[1131],s_t[1131],c_t[1130],c_t2[1131],s_t2[1131]);
fa fau_1_1132(b_i_s[1132],s_t[1132],c_t[1131],c_t2[1132],s_t2[1132]);
fa fau_1_1133(b_i_s[1133],s_t[1133],c_t[1132],c_t2[1133],s_t2[1133]);
fa fau_1_1134(b_i_s[1134],s_t[1134],c_t[1133],c_t2[1134],s_t2[1134]);
fa fau_1_1135(b_i_s[1135],s_t[1135],c_t[1134],c_t2[1135],s_t2[1135]);
fa fau_1_1136(b_i_s[1136],s_t[1136],c_t[1135],c_t2[1136],s_t2[1136]);
fa fau_1_1137(b_i_s[1137],s_t[1137],c_t[1136],c_t2[1137],s_t2[1137]);
fa fau_1_1138(b_i_s[1138],s_t[1138],c_t[1137],c_t2[1138],s_t2[1138]);
fa fau_1_1139(b_i_s[1139],s_t[1139],c_t[1138],c_t2[1139],s_t2[1139]);
fa fau_1_1140(b_i_s[1140],s_t[1140],c_t[1139],c_t2[1140],s_t2[1140]);
fa fau_1_1141(b_i_s[1141],s_t[1141],c_t[1140],c_t2[1141],s_t2[1141]);
fa fau_1_1142(b_i_s[1142],s_t[1142],c_t[1141],c_t2[1142],s_t2[1142]);
fa fau_1_1143(b_i_s[1143],s_t[1143],c_t[1142],c_t2[1143],s_t2[1143]);
fa fau_1_1144(b_i_s[1144],s_t[1144],c_t[1143],c_t2[1144],s_t2[1144]);
fa fau_1_1145(b_i_s[1145],s_t[1145],c_t[1144],c_t2[1145],s_t2[1145]);
fa fau_1_1146(b_i_s[1146],s_t[1146],c_t[1145],c_t2[1146],s_t2[1146]);
fa fau_1_1147(b_i_s[1147],s_t[1147],c_t[1146],c_t2[1147],s_t2[1147]);
fa fau_1_1148(b_i_s[1148],s_t[1148],c_t[1147],c_t2[1148],s_t2[1148]);
fa fau_1_1149(b_i_s[1149],s_t[1149],c_t[1148],c_t2[1149],s_t2[1149]);
fa fau_1_1150(b_i_s[1150],s_t[1150],c_t[1149],c_t2[1150],s_t2[1150]);
fa fau_1_1151(b_i_s[1151],s_t[1151],c_t[1150],c_t2[1151],s_t2[1151]);
fa fau_1_1152(b_i_s[1152],s_t[1152],c_t[1151],c_t2[1152],s_t2[1152]);
fa fau_1_1153(b_i_s[1153],s_t[1153],c_t[1152],c_t2[1153],s_t2[1153]);
fa fau_1_1154(b_i_s[1154],s_t[1154],c_t[1153],c_t2[1154],s_t2[1154]);
fa fau_1_1155(b_i_s[1155],s_t[1155],c_t[1154],c_t2[1155],s_t2[1155]);
fa fau_1_1156(b_i_s[1156],s_t[1156],c_t[1155],c_t2[1156],s_t2[1156]);
fa fau_1_1157(b_i_s[1157],s_t[1157],c_t[1156],c_t2[1157],s_t2[1157]);
fa fau_1_1158(b_i_s[1158],s_t[1158],c_t[1157],c_t2[1158],s_t2[1158]);
fa fau_1_1159(b_i_s[1159],s_t[1159],c_t[1158],c_t2[1159],s_t2[1159]);
fa fau_1_1160(b_i_s[1160],s_t[1160],c_t[1159],c_t2[1160],s_t2[1160]);
fa fau_1_1161(b_i_s[1161],s_t[1161],c_t[1160],c_t2[1161],s_t2[1161]);
fa fau_1_1162(b_i_s[1162],s_t[1162],c_t[1161],c_t2[1162],s_t2[1162]);
fa fau_1_1163(b_i_s[1163],s_t[1163],c_t[1162],c_t2[1163],s_t2[1163]);
fa fau_1_1164(b_i_s[1164],s_t[1164],c_t[1163],c_t2[1164],s_t2[1164]);
fa fau_1_1165(b_i_s[1165],s_t[1165],c_t[1164],c_t2[1165],s_t2[1165]);
fa fau_1_1166(b_i_s[1166],s_t[1166],c_t[1165],c_t2[1166],s_t2[1166]);
fa fau_1_1167(b_i_s[1167],s_t[1167],c_t[1166],c_t2[1167],s_t2[1167]);
fa fau_1_1168(b_i_s[1168],s_t[1168],c_t[1167],c_t2[1168],s_t2[1168]);
fa fau_1_1169(b_i_s[1169],s_t[1169],c_t[1168],c_t2[1169],s_t2[1169]);
fa fau_1_1170(b_i_s[1170],s_t[1170],c_t[1169],c_t2[1170],s_t2[1170]);
fa fau_1_1171(b_i_s[1171],s_t[1171],c_t[1170],c_t2[1171],s_t2[1171]);
fa fau_1_1172(b_i_s[1172],s_t[1172],c_t[1171],c_t2[1172],s_t2[1172]);
fa fau_1_1173(b_i_s[1173],s_t[1173],c_t[1172],c_t2[1173],s_t2[1173]);
fa fau_1_1174(b_i_s[1174],s_t[1174],c_t[1173],c_t2[1174],s_t2[1174]);
fa fau_1_1175(b_i_s[1175],s_t[1175],c_t[1174],c_t2[1175],s_t2[1175]);
fa fau_1_1176(b_i_s[1176],s_t[1176],c_t[1175],c_t2[1176],s_t2[1176]);
fa fau_1_1177(b_i_s[1177],s_t[1177],c_t[1176],c_t2[1177],s_t2[1177]);
fa fau_1_1178(b_i_s[1178],s_t[1178],c_t[1177],c_t2[1178],s_t2[1178]);
fa fau_1_1179(b_i_s[1179],s_t[1179],c_t[1178],c_t2[1179],s_t2[1179]);
fa fau_1_1180(b_i_s[1180],s_t[1180],c_t[1179],c_t2[1180],s_t2[1180]);
fa fau_1_1181(b_i_s[1181],s_t[1181],c_t[1180],c_t2[1181],s_t2[1181]);
fa fau_1_1182(b_i_s[1182],s_t[1182],c_t[1181],c_t2[1182],s_t2[1182]);
fa fau_1_1183(b_i_s[1183],s_t[1183],c_t[1182],c_t2[1183],s_t2[1183]);
fa fau_1_1184(b_i_s[1184],s_t[1184],c_t[1183],c_t2[1184],s_t2[1184]);
fa fau_1_1185(b_i_s[1185],s_t[1185],c_t[1184],c_t2[1185],s_t2[1185]);
fa fau_1_1186(b_i_s[1186],s_t[1186],c_t[1185],c_t2[1186],s_t2[1186]);
fa fau_1_1187(b_i_s[1187],s_t[1187],c_t[1186],c_t2[1187],s_t2[1187]);
fa fau_1_1188(b_i_s[1188],s_t[1188],c_t[1187],c_t2[1188],s_t2[1188]);
fa fau_1_1189(b_i_s[1189],s_t[1189],c_t[1188],c_t2[1189],s_t2[1189]);
fa fau_1_1190(b_i_s[1190],s_t[1190],c_t[1189],c_t2[1190],s_t2[1190]);
fa fau_1_1191(b_i_s[1191],s_t[1191],c_t[1190],c_t2[1191],s_t2[1191]);
fa fau_1_1192(b_i_s[1192],s_t[1192],c_t[1191],c_t2[1192],s_t2[1192]);
fa fau_1_1193(b_i_s[1193],s_t[1193],c_t[1192],c_t2[1193],s_t2[1193]);
fa fau_1_1194(b_i_s[1194],s_t[1194],c_t[1193],c_t2[1194],s_t2[1194]);
fa fau_1_1195(b_i_s[1195],s_t[1195],c_t[1194],c_t2[1195],s_t2[1195]);
fa fau_1_1196(b_i_s[1196],s_t[1196],c_t[1195],c_t2[1196],s_t2[1196]);
fa fau_1_1197(b_i_s[1197],s_t[1197],c_t[1196],c_t2[1197],s_t2[1197]);
fa fau_1_1198(b_i_s[1198],s_t[1198],c_t[1197],c_t2[1198],s_t2[1198]);
fa fau_1_1199(b_i_s[1199],s_t[1199],c_t[1198],c_t2[1199],s_t2[1199]);
fa fau_1_1200(b_i_s[1200],s_t[1200],c_t[1199],c_t2[1200],s_t2[1200]);
fa fau_1_1201(b_i_s[1201],s_t[1201],c_t[1200],c_t2[1201],s_t2[1201]);
fa fau_1_1202(b_i_s[1202],s_t[1202],c_t[1201],c_t2[1202],s_t2[1202]);
fa fau_1_1203(b_i_s[1203],s_t[1203],c_t[1202],c_t2[1203],s_t2[1203]);
fa fau_1_1204(b_i_s[1204],s_t[1204],c_t[1203],c_t2[1204],s_t2[1204]);
fa fau_1_1205(b_i_s[1205],s_t[1205],c_t[1204],c_t2[1205],s_t2[1205]);
fa fau_1_1206(b_i_s[1206],s_t[1206],c_t[1205],c_t2[1206],s_t2[1206]);
fa fau_1_1207(b_i_s[1207],s_t[1207],c_t[1206],c_t2[1207],s_t2[1207]);
fa fau_1_1208(b_i_s[1208],s_t[1208],c_t[1207],c_t2[1208],s_t2[1208]);
fa fau_1_1209(b_i_s[1209],s_t[1209],c_t[1208],c_t2[1209],s_t2[1209]);
fa fau_1_1210(b_i_s[1210],s_t[1210],c_t[1209],c_t2[1210],s_t2[1210]);
fa fau_1_1211(b_i_s[1211],s_t[1211],c_t[1210],c_t2[1211],s_t2[1211]);
fa fau_1_1212(b_i_s[1212],s_t[1212],c_t[1211],c_t2[1212],s_t2[1212]);
fa fau_1_1213(b_i_s[1213],s_t[1213],c_t[1212],c_t2[1213],s_t2[1213]);
fa fau_1_1214(b_i_s[1214],s_t[1214],c_t[1213],c_t2[1214],s_t2[1214]);
fa fau_1_1215(b_i_s[1215],s_t[1215],c_t[1214],c_t2[1215],s_t2[1215]);
fa fau_1_1216(b_i_s[1216],s_t[1216],c_t[1215],c_t2[1216],s_t2[1216]);
fa fau_1_1217(b_i_s[1217],s_t[1217],c_t[1216],c_t2[1217],s_t2[1217]);
fa fau_1_1218(b_i_s[1218],s_t[1218],c_t[1217],c_t2[1218],s_t2[1218]);
fa fau_1_1219(b_i_s[1219],s_t[1219],c_t[1218],c_t2[1219],s_t2[1219]);
fa fau_1_1220(b_i_s[1220],s_t[1220],c_t[1219],c_t2[1220],s_t2[1220]);
fa fau_1_1221(b_i_s[1221],s_t[1221],c_t[1220],c_t2[1221],s_t2[1221]);
fa fau_1_1222(b_i_s[1222],s_t[1222],c_t[1221],c_t2[1222],s_t2[1222]);
fa fau_1_1223(b_i_s[1223],s_t[1223],c_t[1222],c_t2[1223],s_t2[1223]);
fa fau_1_1224(b_i_s[1224],s_t[1224],c_t[1223],c_t2[1224],s_t2[1224]);
fa fau_1_1225(b_i_s[1225],s_t[1225],c_t[1224],c_t2[1225],s_t2[1225]);
fa fau_1_1226(b_i_s[1226],s_t[1226],c_t[1225],c_t2[1226],s_t2[1226]);
fa fau_1_1227(b_i_s[1227],s_t[1227],c_t[1226],c_t2[1227],s_t2[1227]);
fa fau_1_1228(b_i_s[1228],s_t[1228],c_t[1227],c_t2[1228],s_t2[1228]);
fa fau_1_1229(b_i_s[1229],s_t[1229],c_t[1228],c_t2[1229],s_t2[1229]);
fa fau_1_1230(b_i_s[1230],s_t[1230],c_t[1229],c_t2[1230],s_t2[1230]);
fa fau_1_1231(b_i_s[1231],s_t[1231],c_t[1230],c_t2[1231],s_t2[1231]);
fa fau_1_1232(b_i_s[1232],s_t[1232],c_t[1231],c_t2[1232],s_t2[1232]);
fa fau_1_1233(b_i_s[1233],s_t[1233],c_t[1232],c_t2[1233],s_t2[1233]);
fa fau_1_1234(b_i_s[1234],s_t[1234],c_t[1233],c_t2[1234],s_t2[1234]);
fa fau_1_1235(b_i_s[1235],s_t[1235],c_t[1234],c_t2[1235],s_t2[1235]);
fa fau_1_1236(b_i_s[1236],s_t[1236],c_t[1235],c_t2[1236],s_t2[1236]);
fa fau_1_1237(b_i_s[1237],s_t[1237],c_t[1236],c_t2[1237],s_t2[1237]);
fa fau_1_1238(b_i_s[1238],s_t[1238],c_t[1237],c_t2[1238],s_t2[1238]);
fa fau_1_1239(b_i_s[1239],s_t[1239],c_t[1238],c_t2[1239],s_t2[1239]);
fa fau_1_1240(b_i_s[1240],s_t[1240],c_t[1239],c_t2[1240],s_t2[1240]);
fa fau_1_1241(b_i_s[1241],s_t[1241],c_t[1240],c_t2[1241],s_t2[1241]);
fa fau_1_1242(b_i_s[1242],s_t[1242],c_t[1241],c_t2[1242],s_t2[1242]);
fa fau_1_1243(b_i_s[1243],s_t[1243],c_t[1242],c_t2[1243],s_t2[1243]);
fa fau_1_1244(b_i_s[1244],s_t[1244],c_t[1243],c_t2[1244],s_t2[1244]);
fa fau_1_1245(b_i_s[1245],s_t[1245],c_t[1244],c_t2[1245],s_t2[1245]);
fa fau_1_1246(b_i_s[1246],s_t[1246],c_t[1245],c_t2[1246],s_t2[1246]);
fa fau_1_1247(b_i_s[1247],s_t[1247],c_t[1246],c_t2[1247],s_t2[1247]);
fa fau_1_1248(b_i_s[1248],s_t[1248],c_t[1247],c_t2[1248],s_t2[1248]);
fa fau_1_1249(b_i_s[1249],s_t[1249],c_t[1248],c_t2[1249],s_t2[1249]);
fa fau_1_1250(b_i_s[1250],s_t[1250],c_t[1249],c_t2[1250],s_t2[1250]);
fa fau_1_1251(b_i_s[1251],s_t[1251],c_t[1250],c_t2[1251],s_t2[1251]);
fa fau_1_1252(b_i_s[1252],s_t[1252],c_t[1251],c_t2[1252],s_t2[1252]);
fa fau_1_1253(b_i_s[1253],s_t[1253],c_t[1252],c_t2[1253],s_t2[1253]);
fa fau_1_1254(b_i_s[1254],s_t[1254],c_t[1253],c_t2[1254],s_t2[1254]);
fa fau_1_1255(b_i_s[1255],s_t[1255],c_t[1254],c_t2[1255],s_t2[1255]);
fa fau_1_1256(b_i_s[1256],s_t[1256],c_t[1255],c_t2[1256],s_t2[1256]);
fa fau_1_1257(b_i_s[1257],s_t[1257],c_t[1256],c_t2[1257],s_t2[1257]);
fa fau_1_1258(b_i_s[1258],s_t[1258],c_t[1257],c_t2[1258],s_t2[1258]);
fa fau_1_1259(b_i_s[1259],s_t[1259],c_t[1258],c_t2[1259],s_t2[1259]);
fa fau_1_1260(b_i_s[1260],s_t[1260],c_t[1259],c_t2[1260],s_t2[1260]);
fa fau_1_1261(b_i_s[1261],s_t[1261],c_t[1260],c_t2[1261],s_t2[1261]);
fa fau_1_1262(b_i_s[1262],s_t[1262],c_t[1261],c_t2[1262],s_t2[1262]);
fa fau_1_1263(b_i_s[1263],s_t[1263],c_t[1262],c_t2[1263],s_t2[1263]);
fa fau_1_1264(b_i_s[1264],s_t[1264],c_t[1263],c_t2[1264],s_t2[1264]);
fa fau_1_1265(b_i_s[1265],s_t[1265],c_t[1264],c_t2[1265],s_t2[1265]);
fa fau_1_1266(b_i_s[1266],s_t[1266],c_t[1265],c_t2[1266],s_t2[1266]);
fa fau_1_1267(b_i_s[1267],s_t[1267],c_t[1266],c_t2[1267],s_t2[1267]);
fa fau_1_1268(b_i_s[1268],s_t[1268],c_t[1267],c_t2[1268],s_t2[1268]);
fa fau_1_1269(b_i_s[1269],s_t[1269],c_t[1268],c_t2[1269],s_t2[1269]);
fa fau_1_1270(b_i_s[1270],s_t[1270],c_t[1269],c_t2[1270],s_t2[1270]);
fa fau_1_1271(b_i_s[1271],s_t[1271],c_t[1270],c_t2[1271],s_t2[1271]);
fa fau_1_1272(b_i_s[1272],s_t[1272],c_t[1271],c_t2[1272],s_t2[1272]);
fa fau_1_1273(b_i_s[1273],s_t[1273],c_t[1272],c_t2[1273],s_t2[1273]);
fa fau_1_1274(b_i_s[1274],s_t[1274],c_t[1273],c_t2[1274],s_t2[1274]);
fa fau_1_1275(b_i_s[1275],s_t[1275],c_t[1274],c_t2[1275],s_t2[1275]);
fa fau_1_1276(b_i_s[1276],s_t[1276],c_t[1275],c_t2[1276],s_t2[1276]);
fa fau_1_1277(b_i_s[1277],s_t[1277],c_t[1276],c_t2[1277],s_t2[1277]);
fa fau_1_1278(b_i_s[1278],s_t[1278],c_t[1277],c_t2[1278],s_t2[1278]);
fa fau_1_1279(b_i_s[1279],s_t[1279],c_t[1278],c_t2[1279],s_t2[1279]);
fa fau_1_1280(b_i_s[1280],s_t[1280],c_t[1279],c_t2[1280],s_t2[1280]);
fa fau_1_1281(b_i_s[1281],s_t[1281],c_t[1280],c_t2[1281],s_t2[1281]);
fa fau_1_1282(b_i_s[1282],s_t[1282],c_t[1281],c_t2[1282],s_t2[1282]);
fa fau_1_1283(b_i_s[1283],s_t[1283],c_t[1282],c_t2[1283],s_t2[1283]);
fa fau_1_1284(b_i_s[1284],s_t[1284],c_t[1283],c_t2[1284],s_t2[1284]);
fa fau_1_1285(b_i_s[1285],s_t[1285],c_t[1284],c_t2[1285],s_t2[1285]);
fa fau_1_1286(b_i_s[1286],s_t[1286],c_t[1285],c_t2[1286],s_t2[1286]);
fa fau_1_1287(b_i_s[1287],s_t[1287],c_t[1286],c_t2[1287],s_t2[1287]);
fa fau_1_1288(b_i_s[1288],s_t[1288],c_t[1287],c_t2[1288],s_t2[1288]);
fa fau_1_1289(b_i_s[1289],s_t[1289],c_t[1288],c_t2[1289],s_t2[1289]);
fa fau_1_1290(b_i_s[1290],s_t[1290],c_t[1289],c_t2[1290],s_t2[1290]);
fa fau_1_1291(b_i_s[1291],s_t[1291],c_t[1290],c_t2[1291],s_t2[1291]);
fa fau_1_1292(b_i_s[1292],s_t[1292],c_t[1291],c_t2[1292],s_t2[1292]);
fa fau_1_1293(b_i_s[1293],s_t[1293],c_t[1292],c_t2[1293],s_t2[1293]);
fa fau_1_1294(b_i_s[1294],s_t[1294],c_t[1293],c_t2[1294],s_t2[1294]);
fa fau_1_1295(b_i_s[1295],s_t[1295],c_t[1294],c_t2[1295],s_t2[1295]);
fa fau_1_1296(b_i_s[1296],s_t[1296],c_t[1295],c_t2[1296],s_t2[1296]);
fa fau_1_1297(b_i_s[1297],s_t[1297],c_t[1296],c_t2[1297],s_t2[1297]);
fa fau_1_1298(b_i_s[1298],s_t[1298],c_t[1297],c_t2[1298],s_t2[1298]);
fa fau_1_1299(b_i_s[1299],s_t[1299],c_t[1298],c_t2[1299],s_t2[1299]);
fa fau_1_1300(b_i_s[1300],s_t[1300],c_t[1299],c_t2[1300],s_t2[1300]);
fa fau_1_1301(b_i_s[1301],s_t[1301],c_t[1300],c_t2[1301],s_t2[1301]);
fa fau_1_1302(b_i_s[1302],s_t[1302],c_t[1301],c_t2[1302],s_t2[1302]);
fa fau_1_1303(b_i_s[1303],s_t[1303],c_t[1302],c_t2[1303],s_t2[1303]);
fa fau_1_1304(b_i_s[1304],s_t[1304],c_t[1303],c_t2[1304],s_t2[1304]);
fa fau_1_1305(b_i_s[1305],s_t[1305],c_t[1304],c_t2[1305],s_t2[1305]);
fa fau_1_1306(b_i_s[1306],s_t[1306],c_t[1305],c_t2[1306],s_t2[1306]);
fa fau_1_1307(b_i_s[1307],s_t[1307],c_t[1306],c_t2[1307],s_t2[1307]);
fa fau_1_1308(b_i_s[1308],s_t[1308],c_t[1307],c_t2[1308],s_t2[1308]);
fa fau_1_1309(b_i_s[1309],s_t[1309],c_t[1308],c_t2[1309],s_t2[1309]);
fa fau_1_1310(b_i_s[1310],s_t[1310],c_t[1309],c_t2[1310],s_t2[1310]);
fa fau_1_1311(b_i_s[1311],s_t[1311],c_t[1310],c_t2[1311],s_t2[1311]);
fa fau_1_1312(b_i_s[1312],s_t[1312],c_t[1311],c_t2[1312],s_t2[1312]);
fa fau_1_1313(b_i_s[1313],s_t[1313],c_t[1312],c_t2[1313],s_t2[1313]);
fa fau_1_1314(b_i_s[1314],s_t[1314],c_t[1313],c_t2[1314],s_t2[1314]);
fa fau_1_1315(b_i_s[1315],s_t[1315],c_t[1314],c_t2[1315],s_t2[1315]);
fa fau_1_1316(b_i_s[1316],s_t[1316],c_t[1315],c_t2[1316],s_t2[1316]);
fa fau_1_1317(b_i_s[1317],s_t[1317],c_t[1316],c_t2[1317],s_t2[1317]);
fa fau_1_1318(b_i_s[1318],s_t[1318],c_t[1317],c_t2[1318],s_t2[1318]);
fa fau_1_1319(b_i_s[1319],s_t[1319],c_t[1318],c_t2[1319],s_t2[1319]);
fa fau_1_1320(b_i_s[1320],s_t[1320],c_t[1319],c_t2[1320],s_t2[1320]);
fa fau_1_1321(b_i_s[1321],s_t[1321],c_t[1320],c_t2[1321],s_t2[1321]);
fa fau_1_1322(b_i_s[1322],s_t[1322],c_t[1321],c_t2[1322],s_t2[1322]);
fa fau_1_1323(b_i_s[1323],s_t[1323],c_t[1322],c_t2[1323],s_t2[1323]);
fa fau_1_1324(b_i_s[1324],s_t[1324],c_t[1323],c_t2[1324],s_t2[1324]);
fa fau_1_1325(b_i_s[1325],s_t[1325],c_t[1324],c_t2[1325],s_t2[1325]);
fa fau_1_1326(b_i_s[1326],s_t[1326],c_t[1325],c_t2[1326],s_t2[1326]);
fa fau_1_1327(b_i_s[1327],s_t[1327],c_t[1326],c_t2[1327],s_t2[1327]);
fa fau_1_1328(b_i_s[1328],s_t[1328],c_t[1327],c_t2[1328],s_t2[1328]);
fa fau_1_1329(b_i_s[1329],s_t[1329],c_t[1328],c_t2[1329],s_t2[1329]);
fa fau_1_1330(b_i_s[1330],s_t[1330],c_t[1329],c_t2[1330],s_t2[1330]);
fa fau_1_1331(b_i_s[1331],s_t[1331],c_t[1330],c_t2[1331],s_t2[1331]);
fa fau_1_1332(b_i_s[1332],s_t[1332],c_t[1331],c_t2[1332],s_t2[1332]);
fa fau_1_1333(b_i_s[1333],s_t[1333],c_t[1332],c_t2[1333],s_t2[1333]);
fa fau_1_1334(b_i_s[1334],s_t[1334],c_t[1333],c_t2[1334],s_t2[1334]);
fa fau_1_1335(b_i_s[1335],s_t[1335],c_t[1334],c_t2[1335],s_t2[1335]);
fa fau_1_1336(b_i_s[1336],s_t[1336],c_t[1335],c_t2[1336],s_t2[1336]);
fa fau_1_1337(b_i_s[1337],s_t[1337],c_t[1336],c_t2[1337],s_t2[1337]);
fa fau_1_1338(b_i_s[1338],s_t[1338],c_t[1337],c_t2[1338],s_t2[1338]);
fa fau_1_1339(b_i_s[1339],s_t[1339],c_t[1338],c_t2[1339],s_t2[1339]);
fa fau_1_1340(b_i_s[1340],s_t[1340],c_t[1339],c_t2[1340],s_t2[1340]);
fa fau_1_1341(b_i_s[1341],s_t[1341],c_t[1340],c_t2[1341],s_t2[1341]);
fa fau_1_1342(b_i_s[1342],s_t[1342],c_t[1341],c_t2[1342],s_t2[1342]);
fa fau_1_1343(b_i_s[1343],s_t[1343],c_t[1342],c_t2[1343],s_t2[1343]);
fa fau_1_1344(b_i_s[1344],s_t[1344],c_t[1343],c_t2[1344],s_t2[1344]);
fa fau_1_1345(b_i_s[1345],s_t[1345],c_t[1344],c_t2[1345],s_t2[1345]);
fa fau_1_1346(b_i_s[1346],s_t[1346],c_t[1345],c_t2[1346],s_t2[1346]);
fa fau_1_1347(b_i_s[1347],s_t[1347],c_t[1346],c_t2[1347],s_t2[1347]);
fa fau_1_1348(b_i_s[1348],s_t[1348],c_t[1347],c_t2[1348],s_t2[1348]);
fa fau_1_1349(b_i_s[1349],s_t[1349],c_t[1348],c_t2[1349],s_t2[1349]);
fa fau_1_1350(b_i_s[1350],s_t[1350],c_t[1349],c_t2[1350],s_t2[1350]);
fa fau_1_1351(b_i_s[1351],s_t[1351],c_t[1350],c_t2[1351],s_t2[1351]);
fa fau_1_1352(b_i_s[1352],s_t[1352],c_t[1351],c_t2[1352],s_t2[1352]);
fa fau_1_1353(b_i_s[1353],s_t[1353],c_t[1352],c_t2[1353],s_t2[1353]);
fa fau_1_1354(b_i_s[1354],s_t[1354],c_t[1353],c_t2[1354],s_t2[1354]);
fa fau_1_1355(b_i_s[1355],s_t[1355],c_t[1354],c_t2[1355],s_t2[1355]);
fa fau_1_1356(b_i_s[1356],s_t[1356],c_t[1355],c_t2[1356],s_t2[1356]);
fa fau_1_1357(b_i_s[1357],s_t[1357],c_t[1356],c_t2[1357],s_t2[1357]);
fa fau_1_1358(b_i_s[1358],s_t[1358],c_t[1357],c_t2[1358],s_t2[1358]);
fa fau_1_1359(b_i_s[1359],s_t[1359],c_t[1358],c_t2[1359],s_t2[1359]);
fa fau_1_1360(b_i_s[1360],s_t[1360],c_t[1359],c_t2[1360],s_t2[1360]);
fa fau_1_1361(b_i_s[1361],s_t[1361],c_t[1360],c_t2[1361],s_t2[1361]);
fa fau_1_1362(b_i_s[1362],s_t[1362],c_t[1361],c_t2[1362],s_t2[1362]);
fa fau_1_1363(b_i_s[1363],s_t[1363],c_t[1362],c_t2[1363],s_t2[1363]);
fa fau_1_1364(b_i_s[1364],s_t[1364],c_t[1363],c_t2[1364],s_t2[1364]);
fa fau_1_1365(b_i_s[1365],s_t[1365],c_t[1364],c_t2[1365],s_t2[1365]);
fa fau_1_1366(b_i_s[1366],s_t[1366],c_t[1365],c_t2[1366],s_t2[1366]);
fa fau_1_1367(b_i_s[1367],s_t[1367],c_t[1366],c_t2[1367],s_t2[1367]);
fa fau_1_1368(b_i_s[1368],s_t[1368],c_t[1367],c_t2[1368],s_t2[1368]);
fa fau_1_1369(b_i_s[1369],s_t[1369],c_t[1368],c_t2[1369],s_t2[1369]);
fa fau_1_1370(b_i_s[1370],s_t[1370],c_t[1369],c_t2[1370],s_t2[1370]);
fa fau_1_1371(b_i_s[1371],s_t[1371],c_t[1370],c_t2[1371],s_t2[1371]);
fa fau_1_1372(b_i_s[1372],s_t[1372],c_t[1371],c_t2[1372],s_t2[1372]);
fa fau_1_1373(b_i_s[1373],s_t[1373],c_t[1372],c_t2[1373],s_t2[1373]);
fa fau_1_1374(b_i_s[1374],s_t[1374],c_t[1373],c_t2[1374],s_t2[1374]);
fa fau_1_1375(b_i_s[1375],s_t[1375],c_t[1374],c_t2[1375],s_t2[1375]);
fa fau_1_1376(b_i_s[1376],s_t[1376],c_t[1375],c_t2[1376],s_t2[1376]);
fa fau_1_1377(b_i_s[1377],s_t[1377],c_t[1376],c_t2[1377],s_t2[1377]);
fa fau_1_1378(b_i_s[1378],s_t[1378],c_t[1377],c_t2[1378],s_t2[1378]);
fa fau_1_1379(b_i_s[1379],s_t[1379],c_t[1378],c_t2[1379],s_t2[1379]);
fa fau_1_1380(b_i_s[1380],s_t[1380],c_t[1379],c_t2[1380],s_t2[1380]);
fa fau_1_1381(b_i_s[1381],s_t[1381],c_t[1380],c_t2[1381],s_t2[1381]);
fa fau_1_1382(b_i_s[1382],s_t[1382],c_t[1381],c_t2[1382],s_t2[1382]);
fa fau_1_1383(b_i_s[1383],s_t[1383],c_t[1382],c_t2[1383],s_t2[1383]);
fa fau_1_1384(b_i_s[1384],s_t[1384],c_t[1383],c_t2[1384],s_t2[1384]);
fa fau_1_1385(b_i_s[1385],s_t[1385],c_t[1384],c_t2[1385],s_t2[1385]);
fa fau_1_1386(b_i_s[1386],s_t[1386],c_t[1385],c_t2[1386],s_t2[1386]);
fa fau_1_1387(b_i_s[1387],s_t[1387],c_t[1386],c_t2[1387],s_t2[1387]);
fa fau_1_1388(b_i_s[1388],s_t[1388],c_t[1387],c_t2[1388],s_t2[1388]);
fa fau_1_1389(b_i_s[1389],s_t[1389],c_t[1388],c_t2[1389],s_t2[1389]);
fa fau_1_1390(b_i_s[1390],s_t[1390],c_t[1389],c_t2[1390],s_t2[1390]);
fa fau_1_1391(b_i_s[1391],s_t[1391],c_t[1390],c_t2[1391],s_t2[1391]);
fa fau_1_1392(b_i_s[1392],s_t[1392],c_t[1391],c_t2[1392],s_t2[1392]);
fa fau_1_1393(b_i_s[1393],s_t[1393],c_t[1392],c_t2[1393],s_t2[1393]);
fa fau_1_1394(b_i_s[1394],s_t[1394],c_t[1393],c_t2[1394],s_t2[1394]);
fa fau_1_1395(b_i_s[1395],s_t[1395],c_t[1394],c_t2[1395],s_t2[1395]);
fa fau_1_1396(b_i_s[1396],s_t[1396],c_t[1395],c_t2[1396],s_t2[1396]);
fa fau_1_1397(b_i_s[1397],s_t[1397],c_t[1396],c_t2[1397],s_t2[1397]);
fa fau_1_1398(b_i_s[1398],s_t[1398],c_t[1397],c_t2[1398],s_t2[1398]);
fa fau_1_1399(b_i_s[1399],s_t[1399],c_t[1398],c_t2[1399],s_t2[1399]);
fa fau_1_1400(b_i_s[1400],s_t[1400],c_t[1399],c_t2[1400],s_t2[1400]);
fa fau_1_1401(b_i_s[1401],s_t[1401],c_t[1400],c_t2[1401],s_t2[1401]);
fa fau_1_1402(b_i_s[1402],s_t[1402],c_t[1401],c_t2[1402],s_t2[1402]);
fa fau_1_1403(b_i_s[1403],s_t[1403],c_t[1402],c_t2[1403],s_t2[1403]);
fa fau_1_1404(b_i_s[1404],s_t[1404],c_t[1403],c_t2[1404],s_t2[1404]);
fa fau_1_1405(b_i_s[1405],s_t[1405],c_t[1404],c_t2[1405],s_t2[1405]);
fa fau_1_1406(b_i_s[1406],s_t[1406],c_t[1405],c_t2[1406],s_t2[1406]);
fa fau_1_1407(b_i_s[1407],s_t[1407],c_t[1406],c_t2[1407],s_t2[1407]);
fa fau_1_1408(b_i_s[1408],s_t[1408],c_t[1407],c_t2[1408],s_t2[1408]);
fa fau_1_1409(b_i_s[1409],s_t[1409],c_t[1408],c_t2[1409],s_t2[1409]);
fa fau_1_1410(b_i_s[1410],s_t[1410],c_t[1409],c_t2[1410],s_t2[1410]);
fa fau_1_1411(b_i_s[1411],s_t[1411],c_t[1410],c_t2[1411],s_t2[1411]);
fa fau_1_1412(b_i_s[1412],s_t[1412],c_t[1411],c_t2[1412],s_t2[1412]);
fa fau_1_1413(b_i_s[1413],s_t[1413],c_t[1412],c_t2[1413],s_t2[1413]);
fa fau_1_1414(b_i_s[1414],s_t[1414],c_t[1413],c_t2[1414],s_t2[1414]);
fa fau_1_1415(b_i_s[1415],s_t[1415],c_t[1414],c_t2[1415],s_t2[1415]);
fa fau_1_1416(b_i_s[1416],s_t[1416],c_t[1415],c_t2[1416],s_t2[1416]);
fa fau_1_1417(b_i_s[1417],s_t[1417],c_t[1416],c_t2[1417],s_t2[1417]);
fa fau_1_1418(b_i_s[1418],s_t[1418],c_t[1417],c_t2[1418],s_t2[1418]);
fa fau_1_1419(b_i_s[1419],s_t[1419],c_t[1418],c_t2[1419],s_t2[1419]);
fa fau_1_1420(b_i_s[1420],s_t[1420],c_t[1419],c_t2[1420],s_t2[1420]);
fa fau_1_1421(b_i_s[1421],s_t[1421],c_t[1420],c_t2[1421],s_t2[1421]);
fa fau_1_1422(b_i_s[1422],s_t[1422],c_t[1421],c_t2[1422],s_t2[1422]);
fa fau_1_1423(b_i_s[1423],s_t[1423],c_t[1422],c_t2[1423],s_t2[1423]);
fa fau_1_1424(b_i_s[1424],s_t[1424],c_t[1423],c_t2[1424],s_t2[1424]);
fa fau_1_1425(b_i_s[1425],s_t[1425],c_t[1424],c_t2[1425],s_t2[1425]);
fa fau_1_1426(b_i_s[1426],s_t[1426],c_t[1425],c_t2[1426],s_t2[1426]);
fa fau_1_1427(b_i_s[1427],s_t[1427],c_t[1426],c_t2[1427],s_t2[1427]);
fa fau_1_1428(b_i_s[1428],s_t[1428],c_t[1427],c_t2[1428],s_t2[1428]);
fa fau_1_1429(b_i_s[1429],s_t[1429],c_t[1428],c_t2[1429],s_t2[1429]);
fa fau_1_1430(b_i_s[1430],s_t[1430],c_t[1429],c_t2[1430],s_t2[1430]);
fa fau_1_1431(b_i_s[1431],s_t[1431],c_t[1430],c_t2[1431],s_t2[1431]);
fa fau_1_1432(b_i_s[1432],s_t[1432],c_t[1431],c_t2[1432],s_t2[1432]);
fa fau_1_1433(b_i_s[1433],s_t[1433],c_t[1432],c_t2[1433],s_t2[1433]);
fa fau_1_1434(b_i_s[1434],s_t[1434],c_t[1433],c_t2[1434],s_t2[1434]);
fa fau_1_1435(b_i_s[1435],s_t[1435],c_t[1434],c_t2[1435],s_t2[1435]);
fa fau_1_1436(b_i_s[1436],s_t[1436],c_t[1435],c_t2[1436],s_t2[1436]);
fa fau_1_1437(b_i_s[1437],s_t[1437],c_t[1436],c_t2[1437],s_t2[1437]);
fa fau_1_1438(b_i_s[1438],s_t[1438],c_t[1437],c_t2[1438],s_t2[1438]);
fa fau_1_1439(b_i_s[1439],s_t[1439],c_t[1438],c_t2[1439],s_t2[1439]);
fa fau_1_1440(b_i_s[1440],s_t[1440],c_t[1439],c_t2[1440],s_t2[1440]);
fa fau_1_1441(b_i_s[1441],s_t[1441],c_t[1440],c_t2[1441],s_t2[1441]);
fa fau_1_1442(b_i_s[1442],s_t[1442],c_t[1441],c_t2[1442],s_t2[1442]);
fa fau_1_1443(b_i_s[1443],s_t[1443],c_t[1442],c_t2[1443],s_t2[1443]);
fa fau_1_1444(b_i_s[1444],s_t[1444],c_t[1443],c_t2[1444],s_t2[1444]);
fa fau_1_1445(b_i_s[1445],s_t[1445],c_t[1444],c_t2[1445],s_t2[1445]);
fa fau_1_1446(b_i_s[1446],s_t[1446],c_t[1445],c_t2[1446],s_t2[1446]);
fa fau_1_1447(b_i_s[1447],s_t[1447],c_t[1446],c_t2[1447],s_t2[1447]);
fa fau_1_1448(b_i_s[1448],s_t[1448],c_t[1447],c_t2[1448],s_t2[1448]);
fa fau_1_1449(b_i_s[1449],s_t[1449],c_t[1448],c_t2[1449],s_t2[1449]);
fa fau_1_1450(b_i_s[1450],s_t[1450],c_t[1449],c_t2[1450],s_t2[1450]);
fa fau_1_1451(b_i_s[1451],s_t[1451],c_t[1450],c_t2[1451],s_t2[1451]);
fa fau_1_1452(b_i_s[1452],s_t[1452],c_t[1451],c_t2[1452],s_t2[1452]);
fa fau_1_1453(b_i_s[1453],s_t[1453],c_t[1452],c_t2[1453],s_t2[1453]);
fa fau_1_1454(b_i_s[1454],s_t[1454],c_t[1453],c_t2[1454],s_t2[1454]);
fa fau_1_1455(b_i_s[1455],s_t[1455],c_t[1454],c_t2[1455],s_t2[1455]);
fa fau_1_1456(b_i_s[1456],s_t[1456],c_t[1455],c_t2[1456],s_t2[1456]);
fa fau_1_1457(b_i_s[1457],s_t[1457],c_t[1456],c_t2[1457],s_t2[1457]);
fa fau_1_1458(b_i_s[1458],s_t[1458],c_t[1457],c_t2[1458],s_t2[1458]);
fa fau_1_1459(b_i_s[1459],s_t[1459],c_t[1458],c_t2[1459],s_t2[1459]);
fa fau_1_1460(b_i_s[1460],s_t[1460],c_t[1459],c_t2[1460],s_t2[1460]);
fa fau_1_1461(b_i_s[1461],s_t[1461],c_t[1460],c_t2[1461],s_t2[1461]);
fa fau_1_1462(b_i_s[1462],s_t[1462],c_t[1461],c_t2[1462],s_t2[1462]);
fa fau_1_1463(b_i_s[1463],s_t[1463],c_t[1462],c_t2[1463],s_t2[1463]);
fa fau_1_1464(b_i_s[1464],s_t[1464],c_t[1463],c_t2[1464],s_t2[1464]);
fa fau_1_1465(b_i_s[1465],s_t[1465],c_t[1464],c_t2[1465],s_t2[1465]);
fa fau_1_1466(b_i_s[1466],s_t[1466],c_t[1465],c_t2[1466],s_t2[1466]);
fa fau_1_1467(b_i_s[1467],s_t[1467],c_t[1466],c_t2[1467],s_t2[1467]);
fa fau_1_1468(b_i_s[1468],s_t[1468],c_t[1467],c_t2[1468],s_t2[1468]);
fa fau_1_1469(b_i_s[1469],s_t[1469],c_t[1468],c_t2[1469],s_t2[1469]);
fa fau_1_1470(b_i_s[1470],s_t[1470],c_t[1469],c_t2[1470],s_t2[1470]);
fa fau_1_1471(b_i_s[1471],s_t[1471],c_t[1470],c_t2[1471],s_t2[1471]);
fa fau_1_1472(b_i_s[1472],s_t[1472],c_t[1471],c_t2[1472],s_t2[1472]);
fa fau_1_1473(b_i_s[1473],s_t[1473],c_t[1472],c_t2[1473],s_t2[1473]);
fa fau_1_1474(b_i_s[1474],s_t[1474],c_t[1473],c_t2[1474],s_t2[1474]);
fa fau_1_1475(b_i_s[1475],s_t[1475],c_t[1474],c_t2[1475],s_t2[1475]);
fa fau_1_1476(b_i_s[1476],s_t[1476],c_t[1475],c_t2[1476],s_t2[1476]);
fa fau_1_1477(b_i_s[1477],s_t[1477],c_t[1476],c_t2[1477],s_t2[1477]);
fa fau_1_1478(b_i_s[1478],s_t[1478],c_t[1477],c_t2[1478],s_t2[1478]);
fa fau_1_1479(b_i_s[1479],s_t[1479],c_t[1478],c_t2[1479],s_t2[1479]);
fa fau_1_1480(b_i_s[1480],s_t[1480],c_t[1479],c_t2[1480],s_t2[1480]);
fa fau_1_1481(b_i_s[1481],s_t[1481],c_t[1480],c_t2[1481],s_t2[1481]);
fa fau_1_1482(b_i_s[1482],s_t[1482],c_t[1481],c_t2[1482],s_t2[1482]);
fa fau_1_1483(b_i_s[1483],s_t[1483],c_t[1482],c_t2[1483],s_t2[1483]);
fa fau_1_1484(b_i_s[1484],s_t[1484],c_t[1483],c_t2[1484],s_t2[1484]);
fa fau_1_1485(b_i_s[1485],s_t[1485],c_t[1484],c_t2[1485],s_t2[1485]);
fa fau_1_1486(b_i_s[1486],s_t[1486],c_t[1485],c_t2[1486],s_t2[1486]);
fa fau_1_1487(b_i_s[1487],s_t[1487],c_t[1486],c_t2[1487],s_t2[1487]);
fa fau_1_1488(b_i_s[1488],s_t[1488],c_t[1487],c_t2[1488],s_t2[1488]);
fa fau_1_1489(b_i_s[1489],s_t[1489],c_t[1488],c_t2[1489],s_t2[1489]);
fa fau_1_1490(b_i_s[1490],s_t[1490],c_t[1489],c_t2[1490],s_t2[1490]);
fa fau_1_1491(b_i_s[1491],s_t[1491],c_t[1490],c_t2[1491],s_t2[1491]);
fa fau_1_1492(b_i_s[1492],s_t[1492],c_t[1491],c_t2[1492],s_t2[1492]);
fa fau_1_1493(b_i_s[1493],s_t[1493],c_t[1492],c_t2[1493],s_t2[1493]);
fa fau_1_1494(b_i_s[1494],s_t[1494],c_t[1493],c_t2[1494],s_t2[1494]);
fa fau_1_1495(b_i_s[1495],s_t[1495],c_t[1494],c_t2[1495],s_t2[1495]);
fa fau_1_1496(b_i_s[1496],s_t[1496],c_t[1495],c_t2[1496],s_t2[1496]);
fa fau_1_1497(b_i_s[1497],s_t[1497],c_t[1496],c_t2[1497],s_t2[1497]);
fa fau_1_1498(b_i_s[1498],s_t[1498],c_t[1497],c_t2[1498],s_t2[1498]);
fa fau_1_1499(b_i_s[1499],s_t[1499],c_t[1498],c_t2[1499],s_t2[1499]);
fa fau_1_1500(b_i_s[1500],s_t[1500],c_t[1499],c_t2[1500],s_t2[1500]);
fa fau_1_1501(b_i_s[1501],s_t[1501],c_t[1500],c_t2[1501],s_t2[1501]);
fa fau_1_1502(b_i_s[1502],s_t[1502],c_t[1501],c_t2[1502],s_t2[1502]);
fa fau_1_1503(b_i_s[1503],s_t[1503],c_t[1502],c_t2[1503],s_t2[1503]);
fa fau_1_1504(b_i_s[1504],s_t[1504],c_t[1503],c_t2[1504],s_t2[1504]);
fa fau_1_1505(b_i_s[1505],s_t[1505],c_t[1504],c_t2[1505],s_t2[1505]);

fa fau_2(b_i_s[0],s_t[0],1'b0,c_t2[0],s_t2[0]);

assign c = {c_t2,1'b0};
assign s = {c_t[1505],s_t2};

ha ha_red(c[1505],s[1505],ha_c,ha_s);
fa fa_red(c[1506],s[1506],ha_c,fa_c,fa_s);

assign M = {fa_c,fa_s,ha_s};

//LUT for assign corr_add depending on the value of p
add_1506_lut add_1506_lut_i(M,corr_add);

csa_1506 csau({1'b0,c[1504:0]},{1'b0,s[1504:0]},corr_add,c_f,s_f);

assign c_o = c_f;
assign s_o = s_f;

endmodule
    