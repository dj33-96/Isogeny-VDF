
module sub_1506_lut(
    input [3:0] M,
    output reg [1505:0] corr_add
);

always @(*) begin
    case(M)
    4'd0:   corr_add = 1506'h0;
    4'd1:   corr_add = 1506'h20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    4'd2:   corr_add = 1506'h10b6cad46b6070b7ed381d9cea88c74ea092c836403f32b6eb2ac931cabd9bd2a300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
    4'd3:   corr_add = 1506'h16d95a8d6c0e16fda703b39d5118e9d4125906c807e656dd6559263957b37a54600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002;
    4'd4:   corr_add = 1506'h216d95a8d6c0e16fda703b39d5118e9d4125906c807e656dd6559263957b37a54600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002;
    4'd5:   corr_add = 1506'h1224607d42215227c7a858d6bf9a55ebe1b858a2c0bd9824c1805b956038d377e900000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003;
    4'd6:   corr_add = 1506'h2db2b51ad81c2dfb4e07673aa231d3a824b20d900fccadbacab24c72af66f4a8c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004;
    4'd7:   corr_add = 1506'h22db2b51ad81c2dfb4e07673aa231d3a824b20d900fccadbacab24c72af66f4a8c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004;
    4'd8:   corr_add = 1506'h1391f62618e23397a218941094abe48922dde90f413bfd9297d5edf8f5b40b1d2f00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005;
    4'd9:   corr_add = 1506'h448c0fa8442a44f8f50b1ad7f34abd7c370b145817b30498300b72ac071a6efd200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006;
    4'd10:  corr_add = 1506'h2448c0fa8442a44f8f50b1ad7f34abd7c370b145817b30498300b72ac071a6efd200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006;
    4'd11:  corr_add = 1506'h14ff8bceefa315077c88cf4a69bd73266403797bc1ba63006e2b805c8b2f42c27500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007;
    4'd12:  corr_add = 1506'h5b656a35b0385bf69c0ece754463a75049641b201f995b75956498e55ecde951800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008;
    4'd13:  corr_add = 1506'h25b656a35b0385bf69c0ece754463a75049641b201f995b75956498e55ecde951800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008;
    4'd14:  corr_add = 1506'h166d2177c663f67756f90a843ecf01c3a52909e84238c86e448112c020aa7a67bb00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009;
    4'd15:  corr_add = 1506'h723ec4c31c4672f443128212957c91245bbd21e8277fb252fabdbf1eb68163a5e0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a;
    default:corr_add = 0;
    endcase
end

endmodule
    