
module csa_1510 (
    input [1509:0] x,y,z,
    output[1509:0] c,s 
);

wire dummy;

assign c[0] = 1'b0;
    
assign {c[1],s[0]} = (x[0]+y[0]+z[0]);
assign {c[2],s[1]} = (x[1]+y[1]+z[1]);
assign {c[3],s[2]} = (x[2]+y[2]+z[2]);
assign {c[4],s[3]} = (x[3]+y[3]+z[3]);
assign {c[5],s[4]} = (x[4]+y[4]+z[4]);
assign {c[6],s[5]} = (x[5]+y[5]+z[5]);
assign {c[7],s[6]} = (x[6]+y[6]+z[6]);
assign {c[8],s[7]} = (x[7]+y[7]+z[7]);
assign {c[9],s[8]} = (x[8]+y[8]+z[8]);
assign {c[10],s[9]} = (x[9]+y[9]+z[9]);
assign {c[11],s[10]} = (x[10]+y[10]+z[10]);
assign {c[12],s[11]} = (x[11]+y[11]+z[11]);
assign {c[13],s[12]} = (x[12]+y[12]+z[12]);
assign {c[14],s[13]} = (x[13]+y[13]+z[13]);
assign {c[15],s[14]} = (x[14]+y[14]+z[14]);
assign {c[16],s[15]} = (x[15]+y[15]+z[15]);
assign {c[17],s[16]} = (x[16]+y[16]+z[16]);
assign {c[18],s[17]} = (x[17]+y[17]+z[17]);
assign {c[19],s[18]} = (x[18]+y[18]+z[18]);
assign {c[20],s[19]} = (x[19]+y[19]+z[19]);
assign {c[21],s[20]} = (x[20]+y[20]+z[20]);
assign {c[22],s[21]} = (x[21]+y[21]+z[21]);
assign {c[23],s[22]} = (x[22]+y[22]+z[22]);
assign {c[24],s[23]} = (x[23]+y[23]+z[23]);
assign {c[25],s[24]} = (x[24]+y[24]+z[24]);
assign {c[26],s[25]} = (x[25]+y[25]+z[25]);
assign {c[27],s[26]} = (x[26]+y[26]+z[26]);
assign {c[28],s[27]} = (x[27]+y[27]+z[27]);
assign {c[29],s[28]} = (x[28]+y[28]+z[28]);
assign {c[30],s[29]} = (x[29]+y[29]+z[29]);
assign {c[31],s[30]} = (x[30]+y[30]+z[30]);
assign {c[32],s[31]} = (x[31]+y[31]+z[31]);
assign {c[33],s[32]} = (x[32]+y[32]+z[32]);
assign {c[34],s[33]} = (x[33]+y[33]+z[33]);
assign {c[35],s[34]} = (x[34]+y[34]+z[34]);
assign {c[36],s[35]} = (x[35]+y[35]+z[35]);
assign {c[37],s[36]} = (x[36]+y[36]+z[36]);
assign {c[38],s[37]} = (x[37]+y[37]+z[37]);
assign {c[39],s[38]} = (x[38]+y[38]+z[38]);
assign {c[40],s[39]} = (x[39]+y[39]+z[39]);
assign {c[41],s[40]} = (x[40]+y[40]+z[40]);
assign {c[42],s[41]} = (x[41]+y[41]+z[41]);
assign {c[43],s[42]} = (x[42]+y[42]+z[42]);
assign {c[44],s[43]} = (x[43]+y[43]+z[43]);
assign {c[45],s[44]} = (x[44]+y[44]+z[44]);
assign {c[46],s[45]} = (x[45]+y[45]+z[45]);
assign {c[47],s[46]} = (x[46]+y[46]+z[46]);
assign {c[48],s[47]} = (x[47]+y[47]+z[47]);
assign {c[49],s[48]} = (x[48]+y[48]+z[48]);
assign {c[50],s[49]} = (x[49]+y[49]+z[49]);
assign {c[51],s[50]} = (x[50]+y[50]+z[50]);
assign {c[52],s[51]} = (x[51]+y[51]+z[51]);
assign {c[53],s[52]} = (x[52]+y[52]+z[52]);
assign {c[54],s[53]} = (x[53]+y[53]+z[53]);
assign {c[55],s[54]} = (x[54]+y[54]+z[54]);
assign {c[56],s[55]} = (x[55]+y[55]+z[55]);
assign {c[57],s[56]} = (x[56]+y[56]+z[56]);
assign {c[58],s[57]} = (x[57]+y[57]+z[57]);
assign {c[59],s[58]} = (x[58]+y[58]+z[58]);
assign {c[60],s[59]} = (x[59]+y[59]+z[59]);
assign {c[61],s[60]} = (x[60]+y[60]+z[60]);
assign {c[62],s[61]} = (x[61]+y[61]+z[61]);
assign {c[63],s[62]} = (x[62]+y[62]+z[62]);
assign {c[64],s[63]} = (x[63]+y[63]+z[63]);
assign {c[65],s[64]} = (x[64]+y[64]+z[64]);
assign {c[66],s[65]} = (x[65]+y[65]+z[65]);
assign {c[67],s[66]} = (x[66]+y[66]+z[66]);
assign {c[68],s[67]} = (x[67]+y[67]+z[67]);
assign {c[69],s[68]} = (x[68]+y[68]+z[68]);
assign {c[70],s[69]} = (x[69]+y[69]+z[69]);
assign {c[71],s[70]} = (x[70]+y[70]+z[70]);
assign {c[72],s[71]} = (x[71]+y[71]+z[71]);
assign {c[73],s[72]} = (x[72]+y[72]+z[72]);
assign {c[74],s[73]} = (x[73]+y[73]+z[73]);
assign {c[75],s[74]} = (x[74]+y[74]+z[74]);
assign {c[76],s[75]} = (x[75]+y[75]+z[75]);
assign {c[77],s[76]} = (x[76]+y[76]+z[76]);
assign {c[78],s[77]} = (x[77]+y[77]+z[77]);
assign {c[79],s[78]} = (x[78]+y[78]+z[78]);
assign {c[80],s[79]} = (x[79]+y[79]+z[79]);
assign {c[81],s[80]} = (x[80]+y[80]+z[80]);
assign {c[82],s[81]} = (x[81]+y[81]+z[81]);
assign {c[83],s[82]} = (x[82]+y[82]+z[82]);
assign {c[84],s[83]} = (x[83]+y[83]+z[83]);
assign {c[85],s[84]} = (x[84]+y[84]+z[84]);
assign {c[86],s[85]} = (x[85]+y[85]+z[85]);
assign {c[87],s[86]} = (x[86]+y[86]+z[86]);
assign {c[88],s[87]} = (x[87]+y[87]+z[87]);
assign {c[89],s[88]} = (x[88]+y[88]+z[88]);
assign {c[90],s[89]} = (x[89]+y[89]+z[89]);
assign {c[91],s[90]} = (x[90]+y[90]+z[90]);
assign {c[92],s[91]} = (x[91]+y[91]+z[91]);
assign {c[93],s[92]} = (x[92]+y[92]+z[92]);
assign {c[94],s[93]} = (x[93]+y[93]+z[93]);
assign {c[95],s[94]} = (x[94]+y[94]+z[94]);
assign {c[96],s[95]} = (x[95]+y[95]+z[95]);
assign {c[97],s[96]} = (x[96]+y[96]+z[96]);
assign {c[98],s[97]} = (x[97]+y[97]+z[97]);
assign {c[99],s[98]} = (x[98]+y[98]+z[98]);
assign {c[100],s[99]} = (x[99]+y[99]+z[99]);
assign {c[101],s[100]} = (x[100]+y[100]+z[100]);
assign {c[102],s[101]} = (x[101]+y[101]+z[101]);
assign {c[103],s[102]} = (x[102]+y[102]+z[102]);
assign {c[104],s[103]} = (x[103]+y[103]+z[103]);
assign {c[105],s[104]} = (x[104]+y[104]+z[104]);
assign {c[106],s[105]} = (x[105]+y[105]+z[105]);
assign {c[107],s[106]} = (x[106]+y[106]+z[106]);
assign {c[108],s[107]} = (x[107]+y[107]+z[107]);
assign {c[109],s[108]} = (x[108]+y[108]+z[108]);
assign {c[110],s[109]} = (x[109]+y[109]+z[109]);
assign {c[111],s[110]} = (x[110]+y[110]+z[110]);
assign {c[112],s[111]} = (x[111]+y[111]+z[111]);
assign {c[113],s[112]} = (x[112]+y[112]+z[112]);
assign {c[114],s[113]} = (x[113]+y[113]+z[113]);
assign {c[115],s[114]} = (x[114]+y[114]+z[114]);
assign {c[116],s[115]} = (x[115]+y[115]+z[115]);
assign {c[117],s[116]} = (x[116]+y[116]+z[116]);
assign {c[118],s[117]} = (x[117]+y[117]+z[117]);
assign {c[119],s[118]} = (x[118]+y[118]+z[118]);
assign {c[120],s[119]} = (x[119]+y[119]+z[119]);
assign {c[121],s[120]} = (x[120]+y[120]+z[120]);
assign {c[122],s[121]} = (x[121]+y[121]+z[121]);
assign {c[123],s[122]} = (x[122]+y[122]+z[122]);
assign {c[124],s[123]} = (x[123]+y[123]+z[123]);
assign {c[125],s[124]} = (x[124]+y[124]+z[124]);
assign {c[126],s[125]} = (x[125]+y[125]+z[125]);
assign {c[127],s[126]} = (x[126]+y[126]+z[126]);
assign {c[128],s[127]} = (x[127]+y[127]+z[127]);
assign {c[129],s[128]} = (x[128]+y[128]+z[128]);
assign {c[130],s[129]} = (x[129]+y[129]+z[129]);
assign {c[131],s[130]} = (x[130]+y[130]+z[130]);
assign {c[132],s[131]} = (x[131]+y[131]+z[131]);
assign {c[133],s[132]} = (x[132]+y[132]+z[132]);
assign {c[134],s[133]} = (x[133]+y[133]+z[133]);
assign {c[135],s[134]} = (x[134]+y[134]+z[134]);
assign {c[136],s[135]} = (x[135]+y[135]+z[135]);
assign {c[137],s[136]} = (x[136]+y[136]+z[136]);
assign {c[138],s[137]} = (x[137]+y[137]+z[137]);
assign {c[139],s[138]} = (x[138]+y[138]+z[138]);
assign {c[140],s[139]} = (x[139]+y[139]+z[139]);
assign {c[141],s[140]} = (x[140]+y[140]+z[140]);
assign {c[142],s[141]} = (x[141]+y[141]+z[141]);
assign {c[143],s[142]} = (x[142]+y[142]+z[142]);
assign {c[144],s[143]} = (x[143]+y[143]+z[143]);
assign {c[145],s[144]} = (x[144]+y[144]+z[144]);
assign {c[146],s[145]} = (x[145]+y[145]+z[145]);
assign {c[147],s[146]} = (x[146]+y[146]+z[146]);
assign {c[148],s[147]} = (x[147]+y[147]+z[147]);
assign {c[149],s[148]} = (x[148]+y[148]+z[148]);
assign {c[150],s[149]} = (x[149]+y[149]+z[149]);
assign {c[151],s[150]} = (x[150]+y[150]+z[150]);
assign {c[152],s[151]} = (x[151]+y[151]+z[151]);
assign {c[153],s[152]} = (x[152]+y[152]+z[152]);
assign {c[154],s[153]} = (x[153]+y[153]+z[153]);
assign {c[155],s[154]} = (x[154]+y[154]+z[154]);
assign {c[156],s[155]} = (x[155]+y[155]+z[155]);
assign {c[157],s[156]} = (x[156]+y[156]+z[156]);
assign {c[158],s[157]} = (x[157]+y[157]+z[157]);
assign {c[159],s[158]} = (x[158]+y[158]+z[158]);
assign {c[160],s[159]} = (x[159]+y[159]+z[159]);
assign {c[161],s[160]} = (x[160]+y[160]+z[160]);
assign {c[162],s[161]} = (x[161]+y[161]+z[161]);
assign {c[163],s[162]} = (x[162]+y[162]+z[162]);
assign {c[164],s[163]} = (x[163]+y[163]+z[163]);
assign {c[165],s[164]} = (x[164]+y[164]+z[164]);
assign {c[166],s[165]} = (x[165]+y[165]+z[165]);
assign {c[167],s[166]} = (x[166]+y[166]+z[166]);
assign {c[168],s[167]} = (x[167]+y[167]+z[167]);
assign {c[169],s[168]} = (x[168]+y[168]+z[168]);
assign {c[170],s[169]} = (x[169]+y[169]+z[169]);
assign {c[171],s[170]} = (x[170]+y[170]+z[170]);
assign {c[172],s[171]} = (x[171]+y[171]+z[171]);
assign {c[173],s[172]} = (x[172]+y[172]+z[172]);
assign {c[174],s[173]} = (x[173]+y[173]+z[173]);
assign {c[175],s[174]} = (x[174]+y[174]+z[174]);
assign {c[176],s[175]} = (x[175]+y[175]+z[175]);
assign {c[177],s[176]} = (x[176]+y[176]+z[176]);
assign {c[178],s[177]} = (x[177]+y[177]+z[177]);
assign {c[179],s[178]} = (x[178]+y[178]+z[178]);
assign {c[180],s[179]} = (x[179]+y[179]+z[179]);
assign {c[181],s[180]} = (x[180]+y[180]+z[180]);
assign {c[182],s[181]} = (x[181]+y[181]+z[181]);
assign {c[183],s[182]} = (x[182]+y[182]+z[182]);
assign {c[184],s[183]} = (x[183]+y[183]+z[183]);
assign {c[185],s[184]} = (x[184]+y[184]+z[184]);
assign {c[186],s[185]} = (x[185]+y[185]+z[185]);
assign {c[187],s[186]} = (x[186]+y[186]+z[186]);
assign {c[188],s[187]} = (x[187]+y[187]+z[187]);
assign {c[189],s[188]} = (x[188]+y[188]+z[188]);
assign {c[190],s[189]} = (x[189]+y[189]+z[189]);
assign {c[191],s[190]} = (x[190]+y[190]+z[190]);
assign {c[192],s[191]} = (x[191]+y[191]+z[191]);
assign {c[193],s[192]} = (x[192]+y[192]+z[192]);
assign {c[194],s[193]} = (x[193]+y[193]+z[193]);
assign {c[195],s[194]} = (x[194]+y[194]+z[194]);
assign {c[196],s[195]} = (x[195]+y[195]+z[195]);
assign {c[197],s[196]} = (x[196]+y[196]+z[196]);
assign {c[198],s[197]} = (x[197]+y[197]+z[197]);
assign {c[199],s[198]} = (x[198]+y[198]+z[198]);
assign {c[200],s[199]} = (x[199]+y[199]+z[199]);
assign {c[201],s[200]} = (x[200]+y[200]+z[200]);
assign {c[202],s[201]} = (x[201]+y[201]+z[201]);
assign {c[203],s[202]} = (x[202]+y[202]+z[202]);
assign {c[204],s[203]} = (x[203]+y[203]+z[203]);
assign {c[205],s[204]} = (x[204]+y[204]+z[204]);
assign {c[206],s[205]} = (x[205]+y[205]+z[205]);
assign {c[207],s[206]} = (x[206]+y[206]+z[206]);
assign {c[208],s[207]} = (x[207]+y[207]+z[207]);
assign {c[209],s[208]} = (x[208]+y[208]+z[208]);
assign {c[210],s[209]} = (x[209]+y[209]+z[209]);
assign {c[211],s[210]} = (x[210]+y[210]+z[210]);
assign {c[212],s[211]} = (x[211]+y[211]+z[211]);
assign {c[213],s[212]} = (x[212]+y[212]+z[212]);
assign {c[214],s[213]} = (x[213]+y[213]+z[213]);
assign {c[215],s[214]} = (x[214]+y[214]+z[214]);
assign {c[216],s[215]} = (x[215]+y[215]+z[215]);
assign {c[217],s[216]} = (x[216]+y[216]+z[216]);
assign {c[218],s[217]} = (x[217]+y[217]+z[217]);
assign {c[219],s[218]} = (x[218]+y[218]+z[218]);
assign {c[220],s[219]} = (x[219]+y[219]+z[219]);
assign {c[221],s[220]} = (x[220]+y[220]+z[220]);
assign {c[222],s[221]} = (x[221]+y[221]+z[221]);
assign {c[223],s[222]} = (x[222]+y[222]+z[222]);
assign {c[224],s[223]} = (x[223]+y[223]+z[223]);
assign {c[225],s[224]} = (x[224]+y[224]+z[224]);
assign {c[226],s[225]} = (x[225]+y[225]+z[225]);
assign {c[227],s[226]} = (x[226]+y[226]+z[226]);
assign {c[228],s[227]} = (x[227]+y[227]+z[227]);
assign {c[229],s[228]} = (x[228]+y[228]+z[228]);
assign {c[230],s[229]} = (x[229]+y[229]+z[229]);
assign {c[231],s[230]} = (x[230]+y[230]+z[230]);
assign {c[232],s[231]} = (x[231]+y[231]+z[231]);
assign {c[233],s[232]} = (x[232]+y[232]+z[232]);
assign {c[234],s[233]} = (x[233]+y[233]+z[233]);
assign {c[235],s[234]} = (x[234]+y[234]+z[234]);
assign {c[236],s[235]} = (x[235]+y[235]+z[235]);
assign {c[237],s[236]} = (x[236]+y[236]+z[236]);
assign {c[238],s[237]} = (x[237]+y[237]+z[237]);
assign {c[239],s[238]} = (x[238]+y[238]+z[238]);
assign {c[240],s[239]} = (x[239]+y[239]+z[239]);
assign {c[241],s[240]} = (x[240]+y[240]+z[240]);
assign {c[242],s[241]} = (x[241]+y[241]+z[241]);
assign {c[243],s[242]} = (x[242]+y[242]+z[242]);
assign {c[244],s[243]} = (x[243]+y[243]+z[243]);
assign {c[245],s[244]} = (x[244]+y[244]+z[244]);
assign {c[246],s[245]} = (x[245]+y[245]+z[245]);
assign {c[247],s[246]} = (x[246]+y[246]+z[246]);
assign {c[248],s[247]} = (x[247]+y[247]+z[247]);
assign {c[249],s[248]} = (x[248]+y[248]+z[248]);
assign {c[250],s[249]} = (x[249]+y[249]+z[249]);
assign {c[251],s[250]} = (x[250]+y[250]+z[250]);
assign {c[252],s[251]} = (x[251]+y[251]+z[251]);
assign {c[253],s[252]} = (x[252]+y[252]+z[252]);
assign {c[254],s[253]} = (x[253]+y[253]+z[253]);
assign {c[255],s[254]} = (x[254]+y[254]+z[254]);
assign {c[256],s[255]} = (x[255]+y[255]+z[255]);
assign {c[257],s[256]} = (x[256]+y[256]+z[256]);
assign {c[258],s[257]} = (x[257]+y[257]+z[257]);
assign {c[259],s[258]} = (x[258]+y[258]+z[258]);
assign {c[260],s[259]} = (x[259]+y[259]+z[259]);
assign {c[261],s[260]} = (x[260]+y[260]+z[260]);
assign {c[262],s[261]} = (x[261]+y[261]+z[261]);
assign {c[263],s[262]} = (x[262]+y[262]+z[262]);
assign {c[264],s[263]} = (x[263]+y[263]+z[263]);
assign {c[265],s[264]} = (x[264]+y[264]+z[264]);
assign {c[266],s[265]} = (x[265]+y[265]+z[265]);
assign {c[267],s[266]} = (x[266]+y[266]+z[266]);
assign {c[268],s[267]} = (x[267]+y[267]+z[267]);
assign {c[269],s[268]} = (x[268]+y[268]+z[268]);
assign {c[270],s[269]} = (x[269]+y[269]+z[269]);
assign {c[271],s[270]} = (x[270]+y[270]+z[270]);
assign {c[272],s[271]} = (x[271]+y[271]+z[271]);
assign {c[273],s[272]} = (x[272]+y[272]+z[272]);
assign {c[274],s[273]} = (x[273]+y[273]+z[273]);
assign {c[275],s[274]} = (x[274]+y[274]+z[274]);
assign {c[276],s[275]} = (x[275]+y[275]+z[275]);
assign {c[277],s[276]} = (x[276]+y[276]+z[276]);
assign {c[278],s[277]} = (x[277]+y[277]+z[277]);
assign {c[279],s[278]} = (x[278]+y[278]+z[278]);
assign {c[280],s[279]} = (x[279]+y[279]+z[279]);
assign {c[281],s[280]} = (x[280]+y[280]+z[280]);
assign {c[282],s[281]} = (x[281]+y[281]+z[281]);
assign {c[283],s[282]} = (x[282]+y[282]+z[282]);
assign {c[284],s[283]} = (x[283]+y[283]+z[283]);
assign {c[285],s[284]} = (x[284]+y[284]+z[284]);
assign {c[286],s[285]} = (x[285]+y[285]+z[285]);
assign {c[287],s[286]} = (x[286]+y[286]+z[286]);
assign {c[288],s[287]} = (x[287]+y[287]+z[287]);
assign {c[289],s[288]} = (x[288]+y[288]+z[288]);
assign {c[290],s[289]} = (x[289]+y[289]+z[289]);
assign {c[291],s[290]} = (x[290]+y[290]+z[290]);
assign {c[292],s[291]} = (x[291]+y[291]+z[291]);
assign {c[293],s[292]} = (x[292]+y[292]+z[292]);
assign {c[294],s[293]} = (x[293]+y[293]+z[293]);
assign {c[295],s[294]} = (x[294]+y[294]+z[294]);
assign {c[296],s[295]} = (x[295]+y[295]+z[295]);
assign {c[297],s[296]} = (x[296]+y[296]+z[296]);
assign {c[298],s[297]} = (x[297]+y[297]+z[297]);
assign {c[299],s[298]} = (x[298]+y[298]+z[298]);
assign {c[300],s[299]} = (x[299]+y[299]+z[299]);
assign {c[301],s[300]} = (x[300]+y[300]+z[300]);
assign {c[302],s[301]} = (x[301]+y[301]+z[301]);
assign {c[303],s[302]} = (x[302]+y[302]+z[302]);
assign {c[304],s[303]} = (x[303]+y[303]+z[303]);
assign {c[305],s[304]} = (x[304]+y[304]+z[304]);
assign {c[306],s[305]} = (x[305]+y[305]+z[305]);
assign {c[307],s[306]} = (x[306]+y[306]+z[306]);
assign {c[308],s[307]} = (x[307]+y[307]+z[307]);
assign {c[309],s[308]} = (x[308]+y[308]+z[308]);
assign {c[310],s[309]} = (x[309]+y[309]+z[309]);
assign {c[311],s[310]} = (x[310]+y[310]+z[310]);
assign {c[312],s[311]} = (x[311]+y[311]+z[311]);
assign {c[313],s[312]} = (x[312]+y[312]+z[312]);
assign {c[314],s[313]} = (x[313]+y[313]+z[313]);
assign {c[315],s[314]} = (x[314]+y[314]+z[314]);
assign {c[316],s[315]} = (x[315]+y[315]+z[315]);
assign {c[317],s[316]} = (x[316]+y[316]+z[316]);
assign {c[318],s[317]} = (x[317]+y[317]+z[317]);
assign {c[319],s[318]} = (x[318]+y[318]+z[318]);
assign {c[320],s[319]} = (x[319]+y[319]+z[319]);
assign {c[321],s[320]} = (x[320]+y[320]+z[320]);
assign {c[322],s[321]} = (x[321]+y[321]+z[321]);
assign {c[323],s[322]} = (x[322]+y[322]+z[322]);
assign {c[324],s[323]} = (x[323]+y[323]+z[323]);
assign {c[325],s[324]} = (x[324]+y[324]+z[324]);
assign {c[326],s[325]} = (x[325]+y[325]+z[325]);
assign {c[327],s[326]} = (x[326]+y[326]+z[326]);
assign {c[328],s[327]} = (x[327]+y[327]+z[327]);
assign {c[329],s[328]} = (x[328]+y[328]+z[328]);
assign {c[330],s[329]} = (x[329]+y[329]+z[329]);
assign {c[331],s[330]} = (x[330]+y[330]+z[330]);
assign {c[332],s[331]} = (x[331]+y[331]+z[331]);
assign {c[333],s[332]} = (x[332]+y[332]+z[332]);
assign {c[334],s[333]} = (x[333]+y[333]+z[333]);
assign {c[335],s[334]} = (x[334]+y[334]+z[334]);
assign {c[336],s[335]} = (x[335]+y[335]+z[335]);
assign {c[337],s[336]} = (x[336]+y[336]+z[336]);
assign {c[338],s[337]} = (x[337]+y[337]+z[337]);
assign {c[339],s[338]} = (x[338]+y[338]+z[338]);
assign {c[340],s[339]} = (x[339]+y[339]+z[339]);
assign {c[341],s[340]} = (x[340]+y[340]+z[340]);
assign {c[342],s[341]} = (x[341]+y[341]+z[341]);
assign {c[343],s[342]} = (x[342]+y[342]+z[342]);
assign {c[344],s[343]} = (x[343]+y[343]+z[343]);
assign {c[345],s[344]} = (x[344]+y[344]+z[344]);
assign {c[346],s[345]} = (x[345]+y[345]+z[345]);
assign {c[347],s[346]} = (x[346]+y[346]+z[346]);
assign {c[348],s[347]} = (x[347]+y[347]+z[347]);
assign {c[349],s[348]} = (x[348]+y[348]+z[348]);
assign {c[350],s[349]} = (x[349]+y[349]+z[349]);
assign {c[351],s[350]} = (x[350]+y[350]+z[350]);
assign {c[352],s[351]} = (x[351]+y[351]+z[351]);
assign {c[353],s[352]} = (x[352]+y[352]+z[352]);
assign {c[354],s[353]} = (x[353]+y[353]+z[353]);
assign {c[355],s[354]} = (x[354]+y[354]+z[354]);
assign {c[356],s[355]} = (x[355]+y[355]+z[355]);
assign {c[357],s[356]} = (x[356]+y[356]+z[356]);
assign {c[358],s[357]} = (x[357]+y[357]+z[357]);
assign {c[359],s[358]} = (x[358]+y[358]+z[358]);
assign {c[360],s[359]} = (x[359]+y[359]+z[359]);
assign {c[361],s[360]} = (x[360]+y[360]+z[360]);
assign {c[362],s[361]} = (x[361]+y[361]+z[361]);
assign {c[363],s[362]} = (x[362]+y[362]+z[362]);
assign {c[364],s[363]} = (x[363]+y[363]+z[363]);
assign {c[365],s[364]} = (x[364]+y[364]+z[364]);
assign {c[366],s[365]} = (x[365]+y[365]+z[365]);
assign {c[367],s[366]} = (x[366]+y[366]+z[366]);
assign {c[368],s[367]} = (x[367]+y[367]+z[367]);
assign {c[369],s[368]} = (x[368]+y[368]+z[368]);
assign {c[370],s[369]} = (x[369]+y[369]+z[369]);
assign {c[371],s[370]} = (x[370]+y[370]+z[370]);
assign {c[372],s[371]} = (x[371]+y[371]+z[371]);
assign {c[373],s[372]} = (x[372]+y[372]+z[372]);
assign {c[374],s[373]} = (x[373]+y[373]+z[373]);
assign {c[375],s[374]} = (x[374]+y[374]+z[374]);
assign {c[376],s[375]} = (x[375]+y[375]+z[375]);
assign {c[377],s[376]} = (x[376]+y[376]+z[376]);
assign {c[378],s[377]} = (x[377]+y[377]+z[377]);
assign {c[379],s[378]} = (x[378]+y[378]+z[378]);
assign {c[380],s[379]} = (x[379]+y[379]+z[379]);
assign {c[381],s[380]} = (x[380]+y[380]+z[380]);
assign {c[382],s[381]} = (x[381]+y[381]+z[381]);
assign {c[383],s[382]} = (x[382]+y[382]+z[382]);
assign {c[384],s[383]} = (x[383]+y[383]+z[383]);
assign {c[385],s[384]} = (x[384]+y[384]+z[384]);
assign {c[386],s[385]} = (x[385]+y[385]+z[385]);
assign {c[387],s[386]} = (x[386]+y[386]+z[386]);
assign {c[388],s[387]} = (x[387]+y[387]+z[387]);
assign {c[389],s[388]} = (x[388]+y[388]+z[388]);
assign {c[390],s[389]} = (x[389]+y[389]+z[389]);
assign {c[391],s[390]} = (x[390]+y[390]+z[390]);
assign {c[392],s[391]} = (x[391]+y[391]+z[391]);
assign {c[393],s[392]} = (x[392]+y[392]+z[392]);
assign {c[394],s[393]} = (x[393]+y[393]+z[393]);
assign {c[395],s[394]} = (x[394]+y[394]+z[394]);
assign {c[396],s[395]} = (x[395]+y[395]+z[395]);
assign {c[397],s[396]} = (x[396]+y[396]+z[396]);
assign {c[398],s[397]} = (x[397]+y[397]+z[397]);
assign {c[399],s[398]} = (x[398]+y[398]+z[398]);
assign {c[400],s[399]} = (x[399]+y[399]+z[399]);
assign {c[401],s[400]} = (x[400]+y[400]+z[400]);
assign {c[402],s[401]} = (x[401]+y[401]+z[401]);
assign {c[403],s[402]} = (x[402]+y[402]+z[402]);
assign {c[404],s[403]} = (x[403]+y[403]+z[403]);
assign {c[405],s[404]} = (x[404]+y[404]+z[404]);
assign {c[406],s[405]} = (x[405]+y[405]+z[405]);
assign {c[407],s[406]} = (x[406]+y[406]+z[406]);
assign {c[408],s[407]} = (x[407]+y[407]+z[407]);
assign {c[409],s[408]} = (x[408]+y[408]+z[408]);
assign {c[410],s[409]} = (x[409]+y[409]+z[409]);
assign {c[411],s[410]} = (x[410]+y[410]+z[410]);
assign {c[412],s[411]} = (x[411]+y[411]+z[411]);
assign {c[413],s[412]} = (x[412]+y[412]+z[412]);
assign {c[414],s[413]} = (x[413]+y[413]+z[413]);
assign {c[415],s[414]} = (x[414]+y[414]+z[414]);
assign {c[416],s[415]} = (x[415]+y[415]+z[415]);
assign {c[417],s[416]} = (x[416]+y[416]+z[416]);
assign {c[418],s[417]} = (x[417]+y[417]+z[417]);
assign {c[419],s[418]} = (x[418]+y[418]+z[418]);
assign {c[420],s[419]} = (x[419]+y[419]+z[419]);
assign {c[421],s[420]} = (x[420]+y[420]+z[420]);
assign {c[422],s[421]} = (x[421]+y[421]+z[421]);
assign {c[423],s[422]} = (x[422]+y[422]+z[422]);
assign {c[424],s[423]} = (x[423]+y[423]+z[423]);
assign {c[425],s[424]} = (x[424]+y[424]+z[424]);
assign {c[426],s[425]} = (x[425]+y[425]+z[425]);
assign {c[427],s[426]} = (x[426]+y[426]+z[426]);
assign {c[428],s[427]} = (x[427]+y[427]+z[427]);
assign {c[429],s[428]} = (x[428]+y[428]+z[428]);
assign {c[430],s[429]} = (x[429]+y[429]+z[429]);
assign {c[431],s[430]} = (x[430]+y[430]+z[430]);
assign {c[432],s[431]} = (x[431]+y[431]+z[431]);
assign {c[433],s[432]} = (x[432]+y[432]+z[432]);
assign {c[434],s[433]} = (x[433]+y[433]+z[433]);
assign {c[435],s[434]} = (x[434]+y[434]+z[434]);
assign {c[436],s[435]} = (x[435]+y[435]+z[435]);
assign {c[437],s[436]} = (x[436]+y[436]+z[436]);
assign {c[438],s[437]} = (x[437]+y[437]+z[437]);
assign {c[439],s[438]} = (x[438]+y[438]+z[438]);
assign {c[440],s[439]} = (x[439]+y[439]+z[439]);
assign {c[441],s[440]} = (x[440]+y[440]+z[440]);
assign {c[442],s[441]} = (x[441]+y[441]+z[441]);
assign {c[443],s[442]} = (x[442]+y[442]+z[442]);
assign {c[444],s[443]} = (x[443]+y[443]+z[443]);
assign {c[445],s[444]} = (x[444]+y[444]+z[444]);
assign {c[446],s[445]} = (x[445]+y[445]+z[445]);
assign {c[447],s[446]} = (x[446]+y[446]+z[446]);
assign {c[448],s[447]} = (x[447]+y[447]+z[447]);
assign {c[449],s[448]} = (x[448]+y[448]+z[448]);
assign {c[450],s[449]} = (x[449]+y[449]+z[449]);
assign {c[451],s[450]} = (x[450]+y[450]+z[450]);
assign {c[452],s[451]} = (x[451]+y[451]+z[451]);
assign {c[453],s[452]} = (x[452]+y[452]+z[452]);
assign {c[454],s[453]} = (x[453]+y[453]+z[453]);
assign {c[455],s[454]} = (x[454]+y[454]+z[454]);
assign {c[456],s[455]} = (x[455]+y[455]+z[455]);
assign {c[457],s[456]} = (x[456]+y[456]+z[456]);
assign {c[458],s[457]} = (x[457]+y[457]+z[457]);
assign {c[459],s[458]} = (x[458]+y[458]+z[458]);
assign {c[460],s[459]} = (x[459]+y[459]+z[459]);
assign {c[461],s[460]} = (x[460]+y[460]+z[460]);
assign {c[462],s[461]} = (x[461]+y[461]+z[461]);
assign {c[463],s[462]} = (x[462]+y[462]+z[462]);
assign {c[464],s[463]} = (x[463]+y[463]+z[463]);
assign {c[465],s[464]} = (x[464]+y[464]+z[464]);
assign {c[466],s[465]} = (x[465]+y[465]+z[465]);
assign {c[467],s[466]} = (x[466]+y[466]+z[466]);
assign {c[468],s[467]} = (x[467]+y[467]+z[467]);
assign {c[469],s[468]} = (x[468]+y[468]+z[468]);
assign {c[470],s[469]} = (x[469]+y[469]+z[469]);
assign {c[471],s[470]} = (x[470]+y[470]+z[470]);
assign {c[472],s[471]} = (x[471]+y[471]+z[471]);
assign {c[473],s[472]} = (x[472]+y[472]+z[472]);
assign {c[474],s[473]} = (x[473]+y[473]+z[473]);
assign {c[475],s[474]} = (x[474]+y[474]+z[474]);
assign {c[476],s[475]} = (x[475]+y[475]+z[475]);
assign {c[477],s[476]} = (x[476]+y[476]+z[476]);
assign {c[478],s[477]} = (x[477]+y[477]+z[477]);
assign {c[479],s[478]} = (x[478]+y[478]+z[478]);
assign {c[480],s[479]} = (x[479]+y[479]+z[479]);
assign {c[481],s[480]} = (x[480]+y[480]+z[480]);
assign {c[482],s[481]} = (x[481]+y[481]+z[481]);
assign {c[483],s[482]} = (x[482]+y[482]+z[482]);
assign {c[484],s[483]} = (x[483]+y[483]+z[483]);
assign {c[485],s[484]} = (x[484]+y[484]+z[484]);
assign {c[486],s[485]} = (x[485]+y[485]+z[485]);
assign {c[487],s[486]} = (x[486]+y[486]+z[486]);
assign {c[488],s[487]} = (x[487]+y[487]+z[487]);
assign {c[489],s[488]} = (x[488]+y[488]+z[488]);
assign {c[490],s[489]} = (x[489]+y[489]+z[489]);
assign {c[491],s[490]} = (x[490]+y[490]+z[490]);
assign {c[492],s[491]} = (x[491]+y[491]+z[491]);
assign {c[493],s[492]} = (x[492]+y[492]+z[492]);
assign {c[494],s[493]} = (x[493]+y[493]+z[493]);
assign {c[495],s[494]} = (x[494]+y[494]+z[494]);
assign {c[496],s[495]} = (x[495]+y[495]+z[495]);
assign {c[497],s[496]} = (x[496]+y[496]+z[496]);
assign {c[498],s[497]} = (x[497]+y[497]+z[497]);
assign {c[499],s[498]} = (x[498]+y[498]+z[498]);
assign {c[500],s[499]} = (x[499]+y[499]+z[499]);
assign {c[501],s[500]} = (x[500]+y[500]+z[500]);
assign {c[502],s[501]} = (x[501]+y[501]+z[501]);
assign {c[503],s[502]} = (x[502]+y[502]+z[502]);
assign {c[504],s[503]} = (x[503]+y[503]+z[503]);
assign {c[505],s[504]} = (x[504]+y[504]+z[504]);
assign {c[506],s[505]} = (x[505]+y[505]+z[505]);
assign {c[507],s[506]} = (x[506]+y[506]+z[506]);
assign {c[508],s[507]} = (x[507]+y[507]+z[507]);
assign {c[509],s[508]} = (x[508]+y[508]+z[508]);
assign {c[510],s[509]} = (x[509]+y[509]+z[509]);
assign {c[511],s[510]} = (x[510]+y[510]+z[510]);
assign {c[512],s[511]} = (x[511]+y[511]+z[511]);
assign {c[513],s[512]} = (x[512]+y[512]+z[512]);
assign {c[514],s[513]} = (x[513]+y[513]+z[513]);
assign {c[515],s[514]} = (x[514]+y[514]+z[514]);
assign {c[516],s[515]} = (x[515]+y[515]+z[515]);
assign {c[517],s[516]} = (x[516]+y[516]+z[516]);
assign {c[518],s[517]} = (x[517]+y[517]+z[517]);
assign {c[519],s[518]} = (x[518]+y[518]+z[518]);
assign {c[520],s[519]} = (x[519]+y[519]+z[519]);
assign {c[521],s[520]} = (x[520]+y[520]+z[520]);
assign {c[522],s[521]} = (x[521]+y[521]+z[521]);
assign {c[523],s[522]} = (x[522]+y[522]+z[522]);
assign {c[524],s[523]} = (x[523]+y[523]+z[523]);
assign {c[525],s[524]} = (x[524]+y[524]+z[524]);
assign {c[526],s[525]} = (x[525]+y[525]+z[525]);
assign {c[527],s[526]} = (x[526]+y[526]+z[526]);
assign {c[528],s[527]} = (x[527]+y[527]+z[527]);
assign {c[529],s[528]} = (x[528]+y[528]+z[528]);
assign {c[530],s[529]} = (x[529]+y[529]+z[529]);
assign {c[531],s[530]} = (x[530]+y[530]+z[530]);
assign {c[532],s[531]} = (x[531]+y[531]+z[531]);
assign {c[533],s[532]} = (x[532]+y[532]+z[532]);
assign {c[534],s[533]} = (x[533]+y[533]+z[533]);
assign {c[535],s[534]} = (x[534]+y[534]+z[534]);
assign {c[536],s[535]} = (x[535]+y[535]+z[535]);
assign {c[537],s[536]} = (x[536]+y[536]+z[536]);
assign {c[538],s[537]} = (x[537]+y[537]+z[537]);
assign {c[539],s[538]} = (x[538]+y[538]+z[538]);
assign {c[540],s[539]} = (x[539]+y[539]+z[539]);
assign {c[541],s[540]} = (x[540]+y[540]+z[540]);
assign {c[542],s[541]} = (x[541]+y[541]+z[541]);
assign {c[543],s[542]} = (x[542]+y[542]+z[542]);
assign {c[544],s[543]} = (x[543]+y[543]+z[543]);
assign {c[545],s[544]} = (x[544]+y[544]+z[544]);
assign {c[546],s[545]} = (x[545]+y[545]+z[545]);
assign {c[547],s[546]} = (x[546]+y[546]+z[546]);
assign {c[548],s[547]} = (x[547]+y[547]+z[547]);
assign {c[549],s[548]} = (x[548]+y[548]+z[548]);
assign {c[550],s[549]} = (x[549]+y[549]+z[549]);
assign {c[551],s[550]} = (x[550]+y[550]+z[550]);
assign {c[552],s[551]} = (x[551]+y[551]+z[551]);
assign {c[553],s[552]} = (x[552]+y[552]+z[552]);
assign {c[554],s[553]} = (x[553]+y[553]+z[553]);
assign {c[555],s[554]} = (x[554]+y[554]+z[554]);
assign {c[556],s[555]} = (x[555]+y[555]+z[555]);
assign {c[557],s[556]} = (x[556]+y[556]+z[556]);
assign {c[558],s[557]} = (x[557]+y[557]+z[557]);
assign {c[559],s[558]} = (x[558]+y[558]+z[558]);
assign {c[560],s[559]} = (x[559]+y[559]+z[559]);
assign {c[561],s[560]} = (x[560]+y[560]+z[560]);
assign {c[562],s[561]} = (x[561]+y[561]+z[561]);
assign {c[563],s[562]} = (x[562]+y[562]+z[562]);
assign {c[564],s[563]} = (x[563]+y[563]+z[563]);
assign {c[565],s[564]} = (x[564]+y[564]+z[564]);
assign {c[566],s[565]} = (x[565]+y[565]+z[565]);
assign {c[567],s[566]} = (x[566]+y[566]+z[566]);
assign {c[568],s[567]} = (x[567]+y[567]+z[567]);
assign {c[569],s[568]} = (x[568]+y[568]+z[568]);
assign {c[570],s[569]} = (x[569]+y[569]+z[569]);
assign {c[571],s[570]} = (x[570]+y[570]+z[570]);
assign {c[572],s[571]} = (x[571]+y[571]+z[571]);
assign {c[573],s[572]} = (x[572]+y[572]+z[572]);
assign {c[574],s[573]} = (x[573]+y[573]+z[573]);
assign {c[575],s[574]} = (x[574]+y[574]+z[574]);
assign {c[576],s[575]} = (x[575]+y[575]+z[575]);
assign {c[577],s[576]} = (x[576]+y[576]+z[576]);
assign {c[578],s[577]} = (x[577]+y[577]+z[577]);
assign {c[579],s[578]} = (x[578]+y[578]+z[578]);
assign {c[580],s[579]} = (x[579]+y[579]+z[579]);
assign {c[581],s[580]} = (x[580]+y[580]+z[580]);
assign {c[582],s[581]} = (x[581]+y[581]+z[581]);
assign {c[583],s[582]} = (x[582]+y[582]+z[582]);
assign {c[584],s[583]} = (x[583]+y[583]+z[583]);
assign {c[585],s[584]} = (x[584]+y[584]+z[584]);
assign {c[586],s[585]} = (x[585]+y[585]+z[585]);
assign {c[587],s[586]} = (x[586]+y[586]+z[586]);
assign {c[588],s[587]} = (x[587]+y[587]+z[587]);
assign {c[589],s[588]} = (x[588]+y[588]+z[588]);
assign {c[590],s[589]} = (x[589]+y[589]+z[589]);
assign {c[591],s[590]} = (x[590]+y[590]+z[590]);
assign {c[592],s[591]} = (x[591]+y[591]+z[591]);
assign {c[593],s[592]} = (x[592]+y[592]+z[592]);
assign {c[594],s[593]} = (x[593]+y[593]+z[593]);
assign {c[595],s[594]} = (x[594]+y[594]+z[594]);
assign {c[596],s[595]} = (x[595]+y[595]+z[595]);
assign {c[597],s[596]} = (x[596]+y[596]+z[596]);
assign {c[598],s[597]} = (x[597]+y[597]+z[597]);
assign {c[599],s[598]} = (x[598]+y[598]+z[598]);
assign {c[600],s[599]} = (x[599]+y[599]+z[599]);
assign {c[601],s[600]} = (x[600]+y[600]+z[600]);
assign {c[602],s[601]} = (x[601]+y[601]+z[601]);
assign {c[603],s[602]} = (x[602]+y[602]+z[602]);
assign {c[604],s[603]} = (x[603]+y[603]+z[603]);
assign {c[605],s[604]} = (x[604]+y[604]+z[604]);
assign {c[606],s[605]} = (x[605]+y[605]+z[605]);
assign {c[607],s[606]} = (x[606]+y[606]+z[606]);
assign {c[608],s[607]} = (x[607]+y[607]+z[607]);
assign {c[609],s[608]} = (x[608]+y[608]+z[608]);
assign {c[610],s[609]} = (x[609]+y[609]+z[609]);
assign {c[611],s[610]} = (x[610]+y[610]+z[610]);
assign {c[612],s[611]} = (x[611]+y[611]+z[611]);
assign {c[613],s[612]} = (x[612]+y[612]+z[612]);
assign {c[614],s[613]} = (x[613]+y[613]+z[613]);
assign {c[615],s[614]} = (x[614]+y[614]+z[614]);
assign {c[616],s[615]} = (x[615]+y[615]+z[615]);
assign {c[617],s[616]} = (x[616]+y[616]+z[616]);
assign {c[618],s[617]} = (x[617]+y[617]+z[617]);
assign {c[619],s[618]} = (x[618]+y[618]+z[618]);
assign {c[620],s[619]} = (x[619]+y[619]+z[619]);
assign {c[621],s[620]} = (x[620]+y[620]+z[620]);
assign {c[622],s[621]} = (x[621]+y[621]+z[621]);
assign {c[623],s[622]} = (x[622]+y[622]+z[622]);
assign {c[624],s[623]} = (x[623]+y[623]+z[623]);
assign {c[625],s[624]} = (x[624]+y[624]+z[624]);
assign {c[626],s[625]} = (x[625]+y[625]+z[625]);
assign {c[627],s[626]} = (x[626]+y[626]+z[626]);
assign {c[628],s[627]} = (x[627]+y[627]+z[627]);
assign {c[629],s[628]} = (x[628]+y[628]+z[628]);
assign {c[630],s[629]} = (x[629]+y[629]+z[629]);
assign {c[631],s[630]} = (x[630]+y[630]+z[630]);
assign {c[632],s[631]} = (x[631]+y[631]+z[631]);
assign {c[633],s[632]} = (x[632]+y[632]+z[632]);
assign {c[634],s[633]} = (x[633]+y[633]+z[633]);
assign {c[635],s[634]} = (x[634]+y[634]+z[634]);
assign {c[636],s[635]} = (x[635]+y[635]+z[635]);
assign {c[637],s[636]} = (x[636]+y[636]+z[636]);
assign {c[638],s[637]} = (x[637]+y[637]+z[637]);
assign {c[639],s[638]} = (x[638]+y[638]+z[638]);
assign {c[640],s[639]} = (x[639]+y[639]+z[639]);
assign {c[641],s[640]} = (x[640]+y[640]+z[640]);
assign {c[642],s[641]} = (x[641]+y[641]+z[641]);
assign {c[643],s[642]} = (x[642]+y[642]+z[642]);
assign {c[644],s[643]} = (x[643]+y[643]+z[643]);
assign {c[645],s[644]} = (x[644]+y[644]+z[644]);
assign {c[646],s[645]} = (x[645]+y[645]+z[645]);
assign {c[647],s[646]} = (x[646]+y[646]+z[646]);
assign {c[648],s[647]} = (x[647]+y[647]+z[647]);
assign {c[649],s[648]} = (x[648]+y[648]+z[648]);
assign {c[650],s[649]} = (x[649]+y[649]+z[649]);
assign {c[651],s[650]} = (x[650]+y[650]+z[650]);
assign {c[652],s[651]} = (x[651]+y[651]+z[651]);
assign {c[653],s[652]} = (x[652]+y[652]+z[652]);
assign {c[654],s[653]} = (x[653]+y[653]+z[653]);
assign {c[655],s[654]} = (x[654]+y[654]+z[654]);
assign {c[656],s[655]} = (x[655]+y[655]+z[655]);
assign {c[657],s[656]} = (x[656]+y[656]+z[656]);
assign {c[658],s[657]} = (x[657]+y[657]+z[657]);
assign {c[659],s[658]} = (x[658]+y[658]+z[658]);
assign {c[660],s[659]} = (x[659]+y[659]+z[659]);
assign {c[661],s[660]} = (x[660]+y[660]+z[660]);
assign {c[662],s[661]} = (x[661]+y[661]+z[661]);
assign {c[663],s[662]} = (x[662]+y[662]+z[662]);
assign {c[664],s[663]} = (x[663]+y[663]+z[663]);
assign {c[665],s[664]} = (x[664]+y[664]+z[664]);
assign {c[666],s[665]} = (x[665]+y[665]+z[665]);
assign {c[667],s[666]} = (x[666]+y[666]+z[666]);
assign {c[668],s[667]} = (x[667]+y[667]+z[667]);
assign {c[669],s[668]} = (x[668]+y[668]+z[668]);
assign {c[670],s[669]} = (x[669]+y[669]+z[669]);
assign {c[671],s[670]} = (x[670]+y[670]+z[670]);
assign {c[672],s[671]} = (x[671]+y[671]+z[671]);
assign {c[673],s[672]} = (x[672]+y[672]+z[672]);
assign {c[674],s[673]} = (x[673]+y[673]+z[673]);
assign {c[675],s[674]} = (x[674]+y[674]+z[674]);
assign {c[676],s[675]} = (x[675]+y[675]+z[675]);
assign {c[677],s[676]} = (x[676]+y[676]+z[676]);
assign {c[678],s[677]} = (x[677]+y[677]+z[677]);
assign {c[679],s[678]} = (x[678]+y[678]+z[678]);
assign {c[680],s[679]} = (x[679]+y[679]+z[679]);
assign {c[681],s[680]} = (x[680]+y[680]+z[680]);
assign {c[682],s[681]} = (x[681]+y[681]+z[681]);
assign {c[683],s[682]} = (x[682]+y[682]+z[682]);
assign {c[684],s[683]} = (x[683]+y[683]+z[683]);
assign {c[685],s[684]} = (x[684]+y[684]+z[684]);
assign {c[686],s[685]} = (x[685]+y[685]+z[685]);
assign {c[687],s[686]} = (x[686]+y[686]+z[686]);
assign {c[688],s[687]} = (x[687]+y[687]+z[687]);
assign {c[689],s[688]} = (x[688]+y[688]+z[688]);
assign {c[690],s[689]} = (x[689]+y[689]+z[689]);
assign {c[691],s[690]} = (x[690]+y[690]+z[690]);
assign {c[692],s[691]} = (x[691]+y[691]+z[691]);
assign {c[693],s[692]} = (x[692]+y[692]+z[692]);
assign {c[694],s[693]} = (x[693]+y[693]+z[693]);
assign {c[695],s[694]} = (x[694]+y[694]+z[694]);
assign {c[696],s[695]} = (x[695]+y[695]+z[695]);
assign {c[697],s[696]} = (x[696]+y[696]+z[696]);
assign {c[698],s[697]} = (x[697]+y[697]+z[697]);
assign {c[699],s[698]} = (x[698]+y[698]+z[698]);
assign {c[700],s[699]} = (x[699]+y[699]+z[699]);
assign {c[701],s[700]} = (x[700]+y[700]+z[700]);
assign {c[702],s[701]} = (x[701]+y[701]+z[701]);
assign {c[703],s[702]} = (x[702]+y[702]+z[702]);
assign {c[704],s[703]} = (x[703]+y[703]+z[703]);
assign {c[705],s[704]} = (x[704]+y[704]+z[704]);
assign {c[706],s[705]} = (x[705]+y[705]+z[705]);
assign {c[707],s[706]} = (x[706]+y[706]+z[706]);
assign {c[708],s[707]} = (x[707]+y[707]+z[707]);
assign {c[709],s[708]} = (x[708]+y[708]+z[708]);
assign {c[710],s[709]} = (x[709]+y[709]+z[709]);
assign {c[711],s[710]} = (x[710]+y[710]+z[710]);
assign {c[712],s[711]} = (x[711]+y[711]+z[711]);
assign {c[713],s[712]} = (x[712]+y[712]+z[712]);
assign {c[714],s[713]} = (x[713]+y[713]+z[713]);
assign {c[715],s[714]} = (x[714]+y[714]+z[714]);
assign {c[716],s[715]} = (x[715]+y[715]+z[715]);
assign {c[717],s[716]} = (x[716]+y[716]+z[716]);
assign {c[718],s[717]} = (x[717]+y[717]+z[717]);
assign {c[719],s[718]} = (x[718]+y[718]+z[718]);
assign {c[720],s[719]} = (x[719]+y[719]+z[719]);
assign {c[721],s[720]} = (x[720]+y[720]+z[720]);
assign {c[722],s[721]} = (x[721]+y[721]+z[721]);
assign {c[723],s[722]} = (x[722]+y[722]+z[722]);
assign {c[724],s[723]} = (x[723]+y[723]+z[723]);
assign {c[725],s[724]} = (x[724]+y[724]+z[724]);
assign {c[726],s[725]} = (x[725]+y[725]+z[725]);
assign {c[727],s[726]} = (x[726]+y[726]+z[726]);
assign {c[728],s[727]} = (x[727]+y[727]+z[727]);
assign {c[729],s[728]} = (x[728]+y[728]+z[728]);
assign {c[730],s[729]} = (x[729]+y[729]+z[729]);
assign {c[731],s[730]} = (x[730]+y[730]+z[730]);
assign {c[732],s[731]} = (x[731]+y[731]+z[731]);
assign {c[733],s[732]} = (x[732]+y[732]+z[732]);
assign {c[734],s[733]} = (x[733]+y[733]+z[733]);
assign {c[735],s[734]} = (x[734]+y[734]+z[734]);
assign {c[736],s[735]} = (x[735]+y[735]+z[735]);
assign {c[737],s[736]} = (x[736]+y[736]+z[736]);
assign {c[738],s[737]} = (x[737]+y[737]+z[737]);
assign {c[739],s[738]} = (x[738]+y[738]+z[738]);
assign {c[740],s[739]} = (x[739]+y[739]+z[739]);
assign {c[741],s[740]} = (x[740]+y[740]+z[740]);
assign {c[742],s[741]} = (x[741]+y[741]+z[741]);
assign {c[743],s[742]} = (x[742]+y[742]+z[742]);
assign {c[744],s[743]} = (x[743]+y[743]+z[743]);
assign {c[745],s[744]} = (x[744]+y[744]+z[744]);
assign {c[746],s[745]} = (x[745]+y[745]+z[745]);
assign {c[747],s[746]} = (x[746]+y[746]+z[746]);
assign {c[748],s[747]} = (x[747]+y[747]+z[747]);
assign {c[749],s[748]} = (x[748]+y[748]+z[748]);
assign {c[750],s[749]} = (x[749]+y[749]+z[749]);
assign {c[751],s[750]} = (x[750]+y[750]+z[750]);
assign {c[752],s[751]} = (x[751]+y[751]+z[751]);
assign {c[753],s[752]} = (x[752]+y[752]+z[752]);
assign {c[754],s[753]} = (x[753]+y[753]+z[753]);
assign {c[755],s[754]} = (x[754]+y[754]+z[754]);
assign {c[756],s[755]} = (x[755]+y[755]+z[755]);
assign {c[757],s[756]} = (x[756]+y[756]+z[756]);
assign {c[758],s[757]} = (x[757]+y[757]+z[757]);
assign {c[759],s[758]} = (x[758]+y[758]+z[758]);
assign {c[760],s[759]} = (x[759]+y[759]+z[759]);
assign {c[761],s[760]} = (x[760]+y[760]+z[760]);
assign {c[762],s[761]} = (x[761]+y[761]+z[761]);
assign {c[763],s[762]} = (x[762]+y[762]+z[762]);
assign {c[764],s[763]} = (x[763]+y[763]+z[763]);
assign {c[765],s[764]} = (x[764]+y[764]+z[764]);
assign {c[766],s[765]} = (x[765]+y[765]+z[765]);
assign {c[767],s[766]} = (x[766]+y[766]+z[766]);
assign {c[768],s[767]} = (x[767]+y[767]+z[767]);
assign {c[769],s[768]} = (x[768]+y[768]+z[768]);
assign {c[770],s[769]} = (x[769]+y[769]+z[769]);
assign {c[771],s[770]} = (x[770]+y[770]+z[770]);
assign {c[772],s[771]} = (x[771]+y[771]+z[771]);
assign {c[773],s[772]} = (x[772]+y[772]+z[772]);
assign {c[774],s[773]} = (x[773]+y[773]+z[773]);
assign {c[775],s[774]} = (x[774]+y[774]+z[774]);
assign {c[776],s[775]} = (x[775]+y[775]+z[775]);
assign {c[777],s[776]} = (x[776]+y[776]+z[776]);
assign {c[778],s[777]} = (x[777]+y[777]+z[777]);
assign {c[779],s[778]} = (x[778]+y[778]+z[778]);
assign {c[780],s[779]} = (x[779]+y[779]+z[779]);
assign {c[781],s[780]} = (x[780]+y[780]+z[780]);
assign {c[782],s[781]} = (x[781]+y[781]+z[781]);
assign {c[783],s[782]} = (x[782]+y[782]+z[782]);
assign {c[784],s[783]} = (x[783]+y[783]+z[783]);
assign {c[785],s[784]} = (x[784]+y[784]+z[784]);
assign {c[786],s[785]} = (x[785]+y[785]+z[785]);
assign {c[787],s[786]} = (x[786]+y[786]+z[786]);
assign {c[788],s[787]} = (x[787]+y[787]+z[787]);
assign {c[789],s[788]} = (x[788]+y[788]+z[788]);
assign {c[790],s[789]} = (x[789]+y[789]+z[789]);
assign {c[791],s[790]} = (x[790]+y[790]+z[790]);
assign {c[792],s[791]} = (x[791]+y[791]+z[791]);
assign {c[793],s[792]} = (x[792]+y[792]+z[792]);
assign {c[794],s[793]} = (x[793]+y[793]+z[793]);
assign {c[795],s[794]} = (x[794]+y[794]+z[794]);
assign {c[796],s[795]} = (x[795]+y[795]+z[795]);
assign {c[797],s[796]} = (x[796]+y[796]+z[796]);
assign {c[798],s[797]} = (x[797]+y[797]+z[797]);
assign {c[799],s[798]} = (x[798]+y[798]+z[798]);
assign {c[800],s[799]} = (x[799]+y[799]+z[799]);
assign {c[801],s[800]} = (x[800]+y[800]+z[800]);
assign {c[802],s[801]} = (x[801]+y[801]+z[801]);
assign {c[803],s[802]} = (x[802]+y[802]+z[802]);
assign {c[804],s[803]} = (x[803]+y[803]+z[803]);
assign {c[805],s[804]} = (x[804]+y[804]+z[804]);
assign {c[806],s[805]} = (x[805]+y[805]+z[805]);
assign {c[807],s[806]} = (x[806]+y[806]+z[806]);
assign {c[808],s[807]} = (x[807]+y[807]+z[807]);
assign {c[809],s[808]} = (x[808]+y[808]+z[808]);
assign {c[810],s[809]} = (x[809]+y[809]+z[809]);
assign {c[811],s[810]} = (x[810]+y[810]+z[810]);
assign {c[812],s[811]} = (x[811]+y[811]+z[811]);
assign {c[813],s[812]} = (x[812]+y[812]+z[812]);
assign {c[814],s[813]} = (x[813]+y[813]+z[813]);
assign {c[815],s[814]} = (x[814]+y[814]+z[814]);
assign {c[816],s[815]} = (x[815]+y[815]+z[815]);
assign {c[817],s[816]} = (x[816]+y[816]+z[816]);
assign {c[818],s[817]} = (x[817]+y[817]+z[817]);
assign {c[819],s[818]} = (x[818]+y[818]+z[818]);
assign {c[820],s[819]} = (x[819]+y[819]+z[819]);
assign {c[821],s[820]} = (x[820]+y[820]+z[820]);
assign {c[822],s[821]} = (x[821]+y[821]+z[821]);
assign {c[823],s[822]} = (x[822]+y[822]+z[822]);
assign {c[824],s[823]} = (x[823]+y[823]+z[823]);
assign {c[825],s[824]} = (x[824]+y[824]+z[824]);
assign {c[826],s[825]} = (x[825]+y[825]+z[825]);
assign {c[827],s[826]} = (x[826]+y[826]+z[826]);
assign {c[828],s[827]} = (x[827]+y[827]+z[827]);
assign {c[829],s[828]} = (x[828]+y[828]+z[828]);
assign {c[830],s[829]} = (x[829]+y[829]+z[829]);
assign {c[831],s[830]} = (x[830]+y[830]+z[830]);
assign {c[832],s[831]} = (x[831]+y[831]+z[831]);
assign {c[833],s[832]} = (x[832]+y[832]+z[832]);
assign {c[834],s[833]} = (x[833]+y[833]+z[833]);
assign {c[835],s[834]} = (x[834]+y[834]+z[834]);
assign {c[836],s[835]} = (x[835]+y[835]+z[835]);
assign {c[837],s[836]} = (x[836]+y[836]+z[836]);
assign {c[838],s[837]} = (x[837]+y[837]+z[837]);
assign {c[839],s[838]} = (x[838]+y[838]+z[838]);
assign {c[840],s[839]} = (x[839]+y[839]+z[839]);
assign {c[841],s[840]} = (x[840]+y[840]+z[840]);
assign {c[842],s[841]} = (x[841]+y[841]+z[841]);
assign {c[843],s[842]} = (x[842]+y[842]+z[842]);
assign {c[844],s[843]} = (x[843]+y[843]+z[843]);
assign {c[845],s[844]} = (x[844]+y[844]+z[844]);
assign {c[846],s[845]} = (x[845]+y[845]+z[845]);
assign {c[847],s[846]} = (x[846]+y[846]+z[846]);
assign {c[848],s[847]} = (x[847]+y[847]+z[847]);
assign {c[849],s[848]} = (x[848]+y[848]+z[848]);
assign {c[850],s[849]} = (x[849]+y[849]+z[849]);
assign {c[851],s[850]} = (x[850]+y[850]+z[850]);
assign {c[852],s[851]} = (x[851]+y[851]+z[851]);
assign {c[853],s[852]} = (x[852]+y[852]+z[852]);
assign {c[854],s[853]} = (x[853]+y[853]+z[853]);
assign {c[855],s[854]} = (x[854]+y[854]+z[854]);
assign {c[856],s[855]} = (x[855]+y[855]+z[855]);
assign {c[857],s[856]} = (x[856]+y[856]+z[856]);
assign {c[858],s[857]} = (x[857]+y[857]+z[857]);
assign {c[859],s[858]} = (x[858]+y[858]+z[858]);
assign {c[860],s[859]} = (x[859]+y[859]+z[859]);
assign {c[861],s[860]} = (x[860]+y[860]+z[860]);
assign {c[862],s[861]} = (x[861]+y[861]+z[861]);
assign {c[863],s[862]} = (x[862]+y[862]+z[862]);
assign {c[864],s[863]} = (x[863]+y[863]+z[863]);
assign {c[865],s[864]} = (x[864]+y[864]+z[864]);
assign {c[866],s[865]} = (x[865]+y[865]+z[865]);
assign {c[867],s[866]} = (x[866]+y[866]+z[866]);
assign {c[868],s[867]} = (x[867]+y[867]+z[867]);
assign {c[869],s[868]} = (x[868]+y[868]+z[868]);
assign {c[870],s[869]} = (x[869]+y[869]+z[869]);
assign {c[871],s[870]} = (x[870]+y[870]+z[870]);
assign {c[872],s[871]} = (x[871]+y[871]+z[871]);
assign {c[873],s[872]} = (x[872]+y[872]+z[872]);
assign {c[874],s[873]} = (x[873]+y[873]+z[873]);
assign {c[875],s[874]} = (x[874]+y[874]+z[874]);
assign {c[876],s[875]} = (x[875]+y[875]+z[875]);
assign {c[877],s[876]} = (x[876]+y[876]+z[876]);
assign {c[878],s[877]} = (x[877]+y[877]+z[877]);
assign {c[879],s[878]} = (x[878]+y[878]+z[878]);
assign {c[880],s[879]} = (x[879]+y[879]+z[879]);
assign {c[881],s[880]} = (x[880]+y[880]+z[880]);
assign {c[882],s[881]} = (x[881]+y[881]+z[881]);
assign {c[883],s[882]} = (x[882]+y[882]+z[882]);
assign {c[884],s[883]} = (x[883]+y[883]+z[883]);
assign {c[885],s[884]} = (x[884]+y[884]+z[884]);
assign {c[886],s[885]} = (x[885]+y[885]+z[885]);
assign {c[887],s[886]} = (x[886]+y[886]+z[886]);
assign {c[888],s[887]} = (x[887]+y[887]+z[887]);
assign {c[889],s[888]} = (x[888]+y[888]+z[888]);
assign {c[890],s[889]} = (x[889]+y[889]+z[889]);
assign {c[891],s[890]} = (x[890]+y[890]+z[890]);
assign {c[892],s[891]} = (x[891]+y[891]+z[891]);
assign {c[893],s[892]} = (x[892]+y[892]+z[892]);
assign {c[894],s[893]} = (x[893]+y[893]+z[893]);
assign {c[895],s[894]} = (x[894]+y[894]+z[894]);
assign {c[896],s[895]} = (x[895]+y[895]+z[895]);
assign {c[897],s[896]} = (x[896]+y[896]+z[896]);
assign {c[898],s[897]} = (x[897]+y[897]+z[897]);
assign {c[899],s[898]} = (x[898]+y[898]+z[898]);
assign {c[900],s[899]} = (x[899]+y[899]+z[899]);
assign {c[901],s[900]} = (x[900]+y[900]+z[900]);
assign {c[902],s[901]} = (x[901]+y[901]+z[901]);
assign {c[903],s[902]} = (x[902]+y[902]+z[902]);
assign {c[904],s[903]} = (x[903]+y[903]+z[903]);
assign {c[905],s[904]} = (x[904]+y[904]+z[904]);
assign {c[906],s[905]} = (x[905]+y[905]+z[905]);
assign {c[907],s[906]} = (x[906]+y[906]+z[906]);
assign {c[908],s[907]} = (x[907]+y[907]+z[907]);
assign {c[909],s[908]} = (x[908]+y[908]+z[908]);
assign {c[910],s[909]} = (x[909]+y[909]+z[909]);
assign {c[911],s[910]} = (x[910]+y[910]+z[910]);
assign {c[912],s[911]} = (x[911]+y[911]+z[911]);
assign {c[913],s[912]} = (x[912]+y[912]+z[912]);
assign {c[914],s[913]} = (x[913]+y[913]+z[913]);
assign {c[915],s[914]} = (x[914]+y[914]+z[914]);
assign {c[916],s[915]} = (x[915]+y[915]+z[915]);
assign {c[917],s[916]} = (x[916]+y[916]+z[916]);
assign {c[918],s[917]} = (x[917]+y[917]+z[917]);
assign {c[919],s[918]} = (x[918]+y[918]+z[918]);
assign {c[920],s[919]} = (x[919]+y[919]+z[919]);
assign {c[921],s[920]} = (x[920]+y[920]+z[920]);
assign {c[922],s[921]} = (x[921]+y[921]+z[921]);
assign {c[923],s[922]} = (x[922]+y[922]+z[922]);
assign {c[924],s[923]} = (x[923]+y[923]+z[923]);
assign {c[925],s[924]} = (x[924]+y[924]+z[924]);
assign {c[926],s[925]} = (x[925]+y[925]+z[925]);
assign {c[927],s[926]} = (x[926]+y[926]+z[926]);
assign {c[928],s[927]} = (x[927]+y[927]+z[927]);
assign {c[929],s[928]} = (x[928]+y[928]+z[928]);
assign {c[930],s[929]} = (x[929]+y[929]+z[929]);
assign {c[931],s[930]} = (x[930]+y[930]+z[930]);
assign {c[932],s[931]} = (x[931]+y[931]+z[931]);
assign {c[933],s[932]} = (x[932]+y[932]+z[932]);
assign {c[934],s[933]} = (x[933]+y[933]+z[933]);
assign {c[935],s[934]} = (x[934]+y[934]+z[934]);
assign {c[936],s[935]} = (x[935]+y[935]+z[935]);
assign {c[937],s[936]} = (x[936]+y[936]+z[936]);
assign {c[938],s[937]} = (x[937]+y[937]+z[937]);
assign {c[939],s[938]} = (x[938]+y[938]+z[938]);
assign {c[940],s[939]} = (x[939]+y[939]+z[939]);
assign {c[941],s[940]} = (x[940]+y[940]+z[940]);
assign {c[942],s[941]} = (x[941]+y[941]+z[941]);
assign {c[943],s[942]} = (x[942]+y[942]+z[942]);
assign {c[944],s[943]} = (x[943]+y[943]+z[943]);
assign {c[945],s[944]} = (x[944]+y[944]+z[944]);
assign {c[946],s[945]} = (x[945]+y[945]+z[945]);
assign {c[947],s[946]} = (x[946]+y[946]+z[946]);
assign {c[948],s[947]} = (x[947]+y[947]+z[947]);
assign {c[949],s[948]} = (x[948]+y[948]+z[948]);
assign {c[950],s[949]} = (x[949]+y[949]+z[949]);
assign {c[951],s[950]} = (x[950]+y[950]+z[950]);
assign {c[952],s[951]} = (x[951]+y[951]+z[951]);
assign {c[953],s[952]} = (x[952]+y[952]+z[952]);
assign {c[954],s[953]} = (x[953]+y[953]+z[953]);
assign {c[955],s[954]} = (x[954]+y[954]+z[954]);
assign {c[956],s[955]} = (x[955]+y[955]+z[955]);
assign {c[957],s[956]} = (x[956]+y[956]+z[956]);
assign {c[958],s[957]} = (x[957]+y[957]+z[957]);
assign {c[959],s[958]} = (x[958]+y[958]+z[958]);
assign {c[960],s[959]} = (x[959]+y[959]+z[959]);
assign {c[961],s[960]} = (x[960]+y[960]+z[960]);
assign {c[962],s[961]} = (x[961]+y[961]+z[961]);
assign {c[963],s[962]} = (x[962]+y[962]+z[962]);
assign {c[964],s[963]} = (x[963]+y[963]+z[963]);
assign {c[965],s[964]} = (x[964]+y[964]+z[964]);
assign {c[966],s[965]} = (x[965]+y[965]+z[965]);
assign {c[967],s[966]} = (x[966]+y[966]+z[966]);
assign {c[968],s[967]} = (x[967]+y[967]+z[967]);
assign {c[969],s[968]} = (x[968]+y[968]+z[968]);
assign {c[970],s[969]} = (x[969]+y[969]+z[969]);
assign {c[971],s[970]} = (x[970]+y[970]+z[970]);
assign {c[972],s[971]} = (x[971]+y[971]+z[971]);
assign {c[973],s[972]} = (x[972]+y[972]+z[972]);
assign {c[974],s[973]} = (x[973]+y[973]+z[973]);
assign {c[975],s[974]} = (x[974]+y[974]+z[974]);
assign {c[976],s[975]} = (x[975]+y[975]+z[975]);
assign {c[977],s[976]} = (x[976]+y[976]+z[976]);
assign {c[978],s[977]} = (x[977]+y[977]+z[977]);
assign {c[979],s[978]} = (x[978]+y[978]+z[978]);
assign {c[980],s[979]} = (x[979]+y[979]+z[979]);
assign {c[981],s[980]} = (x[980]+y[980]+z[980]);
assign {c[982],s[981]} = (x[981]+y[981]+z[981]);
assign {c[983],s[982]} = (x[982]+y[982]+z[982]);
assign {c[984],s[983]} = (x[983]+y[983]+z[983]);
assign {c[985],s[984]} = (x[984]+y[984]+z[984]);
assign {c[986],s[985]} = (x[985]+y[985]+z[985]);
assign {c[987],s[986]} = (x[986]+y[986]+z[986]);
assign {c[988],s[987]} = (x[987]+y[987]+z[987]);
assign {c[989],s[988]} = (x[988]+y[988]+z[988]);
assign {c[990],s[989]} = (x[989]+y[989]+z[989]);
assign {c[991],s[990]} = (x[990]+y[990]+z[990]);
assign {c[992],s[991]} = (x[991]+y[991]+z[991]);
assign {c[993],s[992]} = (x[992]+y[992]+z[992]);
assign {c[994],s[993]} = (x[993]+y[993]+z[993]);
assign {c[995],s[994]} = (x[994]+y[994]+z[994]);
assign {c[996],s[995]} = (x[995]+y[995]+z[995]);
assign {c[997],s[996]} = (x[996]+y[996]+z[996]);
assign {c[998],s[997]} = (x[997]+y[997]+z[997]);
assign {c[999],s[998]} = (x[998]+y[998]+z[998]);
assign {c[1000],s[999]} = (x[999]+y[999]+z[999]);
assign {c[1001],s[1000]} = (x[1000]+y[1000]+z[1000]);
assign {c[1002],s[1001]} = (x[1001]+y[1001]+z[1001]);
assign {c[1003],s[1002]} = (x[1002]+y[1002]+z[1002]);
assign {c[1004],s[1003]} = (x[1003]+y[1003]+z[1003]);
assign {c[1005],s[1004]} = (x[1004]+y[1004]+z[1004]);
assign {c[1006],s[1005]} = (x[1005]+y[1005]+z[1005]);
assign {c[1007],s[1006]} = (x[1006]+y[1006]+z[1006]);
assign {c[1008],s[1007]} = (x[1007]+y[1007]+z[1007]);
assign {c[1009],s[1008]} = (x[1008]+y[1008]+z[1008]);
assign {c[1010],s[1009]} = (x[1009]+y[1009]+z[1009]);
assign {c[1011],s[1010]} = (x[1010]+y[1010]+z[1010]);
assign {c[1012],s[1011]} = (x[1011]+y[1011]+z[1011]);
assign {c[1013],s[1012]} = (x[1012]+y[1012]+z[1012]);
assign {c[1014],s[1013]} = (x[1013]+y[1013]+z[1013]);
assign {c[1015],s[1014]} = (x[1014]+y[1014]+z[1014]);
assign {c[1016],s[1015]} = (x[1015]+y[1015]+z[1015]);
assign {c[1017],s[1016]} = (x[1016]+y[1016]+z[1016]);
assign {c[1018],s[1017]} = (x[1017]+y[1017]+z[1017]);
assign {c[1019],s[1018]} = (x[1018]+y[1018]+z[1018]);
assign {c[1020],s[1019]} = (x[1019]+y[1019]+z[1019]);
assign {c[1021],s[1020]} = (x[1020]+y[1020]+z[1020]);
assign {c[1022],s[1021]} = (x[1021]+y[1021]+z[1021]);
assign {c[1023],s[1022]} = (x[1022]+y[1022]+z[1022]);
assign {c[1024],s[1023]} = (x[1023]+y[1023]+z[1023]);
assign {c[1025],s[1024]} = (x[1024]+y[1024]+z[1024]);
assign {c[1026],s[1025]} = (x[1025]+y[1025]+z[1025]);
assign {c[1027],s[1026]} = (x[1026]+y[1026]+z[1026]);
assign {c[1028],s[1027]} = (x[1027]+y[1027]+z[1027]);
assign {c[1029],s[1028]} = (x[1028]+y[1028]+z[1028]);
assign {c[1030],s[1029]} = (x[1029]+y[1029]+z[1029]);
assign {c[1031],s[1030]} = (x[1030]+y[1030]+z[1030]);
assign {c[1032],s[1031]} = (x[1031]+y[1031]+z[1031]);
assign {c[1033],s[1032]} = (x[1032]+y[1032]+z[1032]);
assign {c[1034],s[1033]} = (x[1033]+y[1033]+z[1033]);
assign {c[1035],s[1034]} = (x[1034]+y[1034]+z[1034]);
assign {c[1036],s[1035]} = (x[1035]+y[1035]+z[1035]);
assign {c[1037],s[1036]} = (x[1036]+y[1036]+z[1036]);
assign {c[1038],s[1037]} = (x[1037]+y[1037]+z[1037]);
assign {c[1039],s[1038]} = (x[1038]+y[1038]+z[1038]);
assign {c[1040],s[1039]} = (x[1039]+y[1039]+z[1039]);
assign {c[1041],s[1040]} = (x[1040]+y[1040]+z[1040]);
assign {c[1042],s[1041]} = (x[1041]+y[1041]+z[1041]);
assign {c[1043],s[1042]} = (x[1042]+y[1042]+z[1042]);
assign {c[1044],s[1043]} = (x[1043]+y[1043]+z[1043]);
assign {c[1045],s[1044]} = (x[1044]+y[1044]+z[1044]);
assign {c[1046],s[1045]} = (x[1045]+y[1045]+z[1045]);
assign {c[1047],s[1046]} = (x[1046]+y[1046]+z[1046]);
assign {c[1048],s[1047]} = (x[1047]+y[1047]+z[1047]);
assign {c[1049],s[1048]} = (x[1048]+y[1048]+z[1048]);
assign {c[1050],s[1049]} = (x[1049]+y[1049]+z[1049]);
assign {c[1051],s[1050]} = (x[1050]+y[1050]+z[1050]);
assign {c[1052],s[1051]} = (x[1051]+y[1051]+z[1051]);
assign {c[1053],s[1052]} = (x[1052]+y[1052]+z[1052]);
assign {c[1054],s[1053]} = (x[1053]+y[1053]+z[1053]);
assign {c[1055],s[1054]} = (x[1054]+y[1054]+z[1054]);
assign {c[1056],s[1055]} = (x[1055]+y[1055]+z[1055]);
assign {c[1057],s[1056]} = (x[1056]+y[1056]+z[1056]);
assign {c[1058],s[1057]} = (x[1057]+y[1057]+z[1057]);
assign {c[1059],s[1058]} = (x[1058]+y[1058]+z[1058]);
assign {c[1060],s[1059]} = (x[1059]+y[1059]+z[1059]);
assign {c[1061],s[1060]} = (x[1060]+y[1060]+z[1060]);
assign {c[1062],s[1061]} = (x[1061]+y[1061]+z[1061]);
assign {c[1063],s[1062]} = (x[1062]+y[1062]+z[1062]);
assign {c[1064],s[1063]} = (x[1063]+y[1063]+z[1063]);
assign {c[1065],s[1064]} = (x[1064]+y[1064]+z[1064]);
assign {c[1066],s[1065]} = (x[1065]+y[1065]+z[1065]);
assign {c[1067],s[1066]} = (x[1066]+y[1066]+z[1066]);
assign {c[1068],s[1067]} = (x[1067]+y[1067]+z[1067]);
assign {c[1069],s[1068]} = (x[1068]+y[1068]+z[1068]);
assign {c[1070],s[1069]} = (x[1069]+y[1069]+z[1069]);
assign {c[1071],s[1070]} = (x[1070]+y[1070]+z[1070]);
assign {c[1072],s[1071]} = (x[1071]+y[1071]+z[1071]);
assign {c[1073],s[1072]} = (x[1072]+y[1072]+z[1072]);
assign {c[1074],s[1073]} = (x[1073]+y[1073]+z[1073]);
assign {c[1075],s[1074]} = (x[1074]+y[1074]+z[1074]);
assign {c[1076],s[1075]} = (x[1075]+y[1075]+z[1075]);
assign {c[1077],s[1076]} = (x[1076]+y[1076]+z[1076]);
assign {c[1078],s[1077]} = (x[1077]+y[1077]+z[1077]);
assign {c[1079],s[1078]} = (x[1078]+y[1078]+z[1078]);
assign {c[1080],s[1079]} = (x[1079]+y[1079]+z[1079]);
assign {c[1081],s[1080]} = (x[1080]+y[1080]+z[1080]);
assign {c[1082],s[1081]} = (x[1081]+y[1081]+z[1081]);
assign {c[1083],s[1082]} = (x[1082]+y[1082]+z[1082]);
assign {c[1084],s[1083]} = (x[1083]+y[1083]+z[1083]);
assign {c[1085],s[1084]} = (x[1084]+y[1084]+z[1084]);
assign {c[1086],s[1085]} = (x[1085]+y[1085]+z[1085]);
assign {c[1087],s[1086]} = (x[1086]+y[1086]+z[1086]);
assign {c[1088],s[1087]} = (x[1087]+y[1087]+z[1087]);
assign {c[1089],s[1088]} = (x[1088]+y[1088]+z[1088]);
assign {c[1090],s[1089]} = (x[1089]+y[1089]+z[1089]);
assign {c[1091],s[1090]} = (x[1090]+y[1090]+z[1090]);
assign {c[1092],s[1091]} = (x[1091]+y[1091]+z[1091]);
assign {c[1093],s[1092]} = (x[1092]+y[1092]+z[1092]);
assign {c[1094],s[1093]} = (x[1093]+y[1093]+z[1093]);
assign {c[1095],s[1094]} = (x[1094]+y[1094]+z[1094]);
assign {c[1096],s[1095]} = (x[1095]+y[1095]+z[1095]);
assign {c[1097],s[1096]} = (x[1096]+y[1096]+z[1096]);
assign {c[1098],s[1097]} = (x[1097]+y[1097]+z[1097]);
assign {c[1099],s[1098]} = (x[1098]+y[1098]+z[1098]);
assign {c[1100],s[1099]} = (x[1099]+y[1099]+z[1099]);
assign {c[1101],s[1100]} = (x[1100]+y[1100]+z[1100]);
assign {c[1102],s[1101]} = (x[1101]+y[1101]+z[1101]);
assign {c[1103],s[1102]} = (x[1102]+y[1102]+z[1102]);
assign {c[1104],s[1103]} = (x[1103]+y[1103]+z[1103]);
assign {c[1105],s[1104]} = (x[1104]+y[1104]+z[1104]);
assign {c[1106],s[1105]} = (x[1105]+y[1105]+z[1105]);
assign {c[1107],s[1106]} = (x[1106]+y[1106]+z[1106]);
assign {c[1108],s[1107]} = (x[1107]+y[1107]+z[1107]);
assign {c[1109],s[1108]} = (x[1108]+y[1108]+z[1108]);
assign {c[1110],s[1109]} = (x[1109]+y[1109]+z[1109]);
assign {c[1111],s[1110]} = (x[1110]+y[1110]+z[1110]);
assign {c[1112],s[1111]} = (x[1111]+y[1111]+z[1111]);
assign {c[1113],s[1112]} = (x[1112]+y[1112]+z[1112]);
assign {c[1114],s[1113]} = (x[1113]+y[1113]+z[1113]);
assign {c[1115],s[1114]} = (x[1114]+y[1114]+z[1114]);
assign {c[1116],s[1115]} = (x[1115]+y[1115]+z[1115]);
assign {c[1117],s[1116]} = (x[1116]+y[1116]+z[1116]);
assign {c[1118],s[1117]} = (x[1117]+y[1117]+z[1117]);
assign {c[1119],s[1118]} = (x[1118]+y[1118]+z[1118]);
assign {c[1120],s[1119]} = (x[1119]+y[1119]+z[1119]);
assign {c[1121],s[1120]} = (x[1120]+y[1120]+z[1120]);
assign {c[1122],s[1121]} = (x[1121]+y[1121]+z[1121]);
assign {c[1123],s[1122]} = (x[1122]+y[1122]+z[1122]);
assign {c[1124],s[1123]} = (x[1123]+y[1123]+z[1123]);
assign {c[1125],s[1124]} = (x[1124]+y[1124]+z[1124]);
assign {c[1126],s[1125]} = (x[1125]+y[1125]+z[1125]);
assign {c[1127],s[1126]} = (x[1126]+y[1126]+z[1126]);
assign {c[1128],s[1127]} = (x[1127]+y[1127]+z[1127]);
assign {c[1129],s[1128]} = (x[1128]+y[1128]+z[1128]);
assign {c[1130],s[1129]} = (x[1129]+y[1129]+z[1129]);
assign {c[1131],s[1130]} = (x[1130]+y[1130]+z[1130]);
assign {c[1132],s[1131]} = (x[1131]+y[1131]+z[1131]);
assign {c[1133],s[1132]} = (x[1132]+y[1132]+z[1132]);
assign {c[1134],s[1133]} = (x[1133]+y[1133]+z[1133]);
assign {c[1135],s[1134]} = (x[1134]+y[1134]+z[1134]);
assign {c[1136],s[1135]} = (x[1135]+y[1135]+z[1135]);
assign {c[1137],s[1136]} = (x[1136]+y[1136]+z[1136]);
assign {c[1138],s[1137]} = (x[1137]+y[1137]+z[1137]);
assign {c[1139],s[1138]} = (x[1138]+y[1138]+z[1138]);
assign {c[1140],s[1139]} = (x[1139]+y[1139]+z[1139]);
assign {c[1141],s[1140]} = (x[1140]+y[1140]+z[1140]);
assign {c[1142],s[1141]} = (x[1141]+y[1141]+z[1141]);
assign {c[1143],s[1142]} = (x[1142]+y[1142]+z[1142]);
assign {c[1144],s[1143]} = (x[1143]+y[1143]+z[1143]);
assign {c[1145],s[1144]} = (x[1144]+y[1144]+z[1144]);
assign {c[1146],s[1145]} = (x[1145]+y[1145]+z[1145]);
assign {c[1147],s[1146]} = (x[1146]+y[1146]+z[1146]);
assign {c[1148],s[1147]} = (x[1147]+y[1147]+z[1147]);
assign {c[1149],s[1148]} = (x[1148]+y[1148]+z[1148]);
assign {c[1150],s[1149]} = (x[1149]+y[1149]+z[1149]);
assign {c[1151],s[1150]} = (x[1150]+y[1150]+z[1150]);
assign {c[1152],s[1151]} = (x[1151]+y[1151]+z[1151]);
assign {c[1153],s[1152]} = (x[1152]+y[1152]+z[1152]);
assign {c[1154],s[1153]} = (x[1153]+y[1153]+z[1153]);
assign {c[1155],s[1154]} = (x[1154]+y[1154]+z[1154]);
assign {c[1156],s[1155]} = (x[1155]+y[1155]+z[1155]);
assign {c[1157],s[1156]} = (x[1156]+y[1156]+z[1156]);
assign {c[1158],s[1157]} = (x[1157]+y[1157]+z[1157]);
assign {c[1159],s[1158]} = (x[1158]+y[1158]+z[1158]);
assign {c[1160],s[1159]} = (x[1159]+y[1159]+z[1159]);
assign {c[1161],s[1160]} = (x[1160]+y[1160]+z[1160]);
assign {c[1162],s[1161]} = (x[1161]+y[1161]+z[1161]);
assign {c[1163],s[1162]} = (x[1162]+y[1162]+z[1162]);
assign {c[1164],s[1163]} = (x[1163]+y[1163]+z[1163]);
assign {c[1165],s[1164]} = (x[1164]+y[1164]+z[1164]);
assign {c[1166],s[1165]} = (x[1165]+y[1165]+z[1165]);
assign {c[1167],s[1166]} = (x[1166]+y[1166]+z[1166]);
assign {c[1168],s[1167]} = (x[1167]+y[1167]+z[1167]);
assign {c[1169],s[1168]} = (x[1168]+y[1168]+z[1168]);
assign {c[1170],s[1169]} = (x[1169]+y[1169]+z[1169]);
assign {c[1171],s[1170]} = (x[1170]+y[1170]+z[1170]);
assign {c[1172],s[1171]} = (x[1171]+y[1171]+z[1171]);
assign {c[1173],s[1172]} = (x[1172]+y[1172]+z[1172]);
assign {c[1174],s[1173]} = (x[1173]+y[1173]+z[1173]);
assign {c[1175],s[1174]} = (x[1174]+y[1174]+z[1174]);
assign {c[1176],s[1175]} = (x[1175]+y[1175]+z[1175]);
assign {c[1177],s[1176]} = (x[1176]+y[1176]+z[1176]);
assign {c[1178],s[1177]} = (x[1177]+y[1177]+z[1177]);
assign {c[1179],s[1178]} = (x[1178]+y[1178]+z[1178]);
assign {c[1180],s[1179]} = (x[1179]+y[1179]+z[1179]);
assign {c[1181],s[1180]} = (x[1180]+y[1180]+z[1180]);
assign {c[1182],s[1181]} = (x[1181]+y[1181]+z[1181]);
assign {c[1183],s[1182]} = (x[1182]+y[1182]+z[1182]);
assign {c[1184],s[1183]} = (x[1183]+y[1183]+z[1183]);
assign {c[1185],s[1184]} = (x[1184]+y[1184]+z[1184]);
assign {c[1186],s[1185]} = (x[1185]+y[1185]+z[1185]);
assign {c[1187],s[1186]} = (x[1186]+y[1186]+z[1186]);
assign {c[1188],s[1187]} = (x[1187]+y[1187]+z[1187]);
assign {c[1189],s[1188]} = (x[1188]+y[1188]+z[1188]);
assign {c[1190],s[1189]} = (x[1189]+y[1189]+z[1189]);
assign {c[1191],s[1190]} = (x[1190]+y[1190]+z[1190]);
assign {c[1192],s[1191]} = (x[1191]+y[1191]+z[1191]);
assign {c[1193],s[1192]} = (x[1192]+y[1192]+z[1192]);
assign {c[1194],s[1193]} = (x[1193]+y[1193]+z[1193]);
assign {c[1195],s[1194]} = (x[1194]+y[1194]+z[1194]);
assign {c[1196],s[1195]} = (x[1195]+y[1195]+z[1195]);
assign {c[1197],s[1196]} = (x[1196]+y[1196]+z[1196]);
assign {c[1198],s[1197]} = (x[1197]+y[1197]+z[1197]);
assign {c[1199],s[1198]} = (x[1198]+y[1198]+z[1198]);
assign {c[1200],s[1199]} = (x[1199]+y[1199]+z[1199]);
assign {c[1201],s[1200]} = (x[1200]+y[1200]+z[1200]);
assign {c[1202],s[1201]} = (x[1201]+y[1201]+z[1201]);
assign {c[1203],s[1202]} = (x[1202]+y[1202]+z[1202]);
assign {c[1204],s[1203]} = (x[1203]+y[1203]+z[1203]);
assign {c[1205],s[1204]} = (x[1204]+y[1204]+z[1204]);
assign {c[1206],s[1205]} = (x[1205]+y[1205]+z[1205]);
assign {c[1207],s[1206]} = (x[1206]+y[1206]+z[1206]);
assign {c[1208],s[1207]} = (x[1207]+y[1207]+z[1207]);
assign {c[1209],s[1208]} = (x[1208]+y[1208]+z[1208]);
assign {c[1210],s[1209]} = (x[1209]+y[1209]+z[1209]);
assign {c[1211],s[1210]} = (x[1210]+y[1210]+z[1210]);
assign {c[1212],s[1211]} = (x[1211]+y[1211]+z[1211]);
assign {c[1213],s[1212]} = (x[1212]+y[1212]+z[1212]);
assign {c[1214],s[1213]} = (x[1213]+y[1213]+z[1213]);
assign {c[1215],s[1214]} = (x[1214]+y[1214]+z[1214]);
assign {c[1216],s[1215]} = (x[1215]+y[1215]+z[1215]);
assign {c[1217],s[1216]} = (x[1216]+y[1216]+z[1216]);
assign {c[1218],s[1217]} = (x[1217]+y[1217]+z[1217]);
assign {c[1219],s[1218]} = (x[1218]+y[1218]+z[1218]);
assign {c[1220],s[1219]} = (x[1219]+y[1219]+z[1219]);
assign {c[1221],s[1220]} = (x[1220]+y[1220]+z[1220]);
assign {c[1222],s[1221]} = (x[1221]+y[1221]+z[1221]);
assign {c[1223],s[1222]} = (x[1222]+y[1222]+z[1222]);
assign {c[1224],s[1223]} = (x[1223]+y[1223]+z[1223]);
assign {c[1225],s[1224]} = (x[1224]+y[1224]+z[1224]);
assign {c[1226],s[1225]} = (x[1225]+y[1225]+z[1225]);
assign {c[1227],s[1226]} = (x[1226]+y[1226]+z[1226]);
assign {c[1228],s[1227]} = (x[1227]+y[1227]+z[1227]);
assign {c[1229],s[1228]} = (x[1228]+y[1228]+z[1228]);
assign {c[1230],s[1229]} = (x[1229]+y[1229]+z[1229]);
assign {c[1231],s[1230]} = (x[1230]+y[1230]+z[1230]);
assign {c[1232],s[1231]} = (x[1231]+y[1231]+z[1231]);
assign {c[1233],s[1232]} = (x[1232]+y[1232]+z[1232]);
assign {c[1234],s[1233]} = (x[1233]+y[1233]+z[1233]);
assign {c[1235],s[1234]} = (x[1234]+y[1234]+z[1234]);
assign {c[1236],s[1235]} = (x[1235]+y[1235]+z[1235]);
assign {c[1237],s[1236]} = (x[1236]+y[1236]+z[1236]);
assign {c[1238],s[1237]} = (x[1237]+y[1237]+z[1237]);
assign {c[1239],s[1238]} = (x[1238]+y[1238]+z[1238]);
assign {c[1240],s[1239]} = (x[1239]+y[1239]+z[1239]);
assign {c[1241],s[1240]} = (x[1240]+y[1240]+z[1240]);
assign {c[1242],s[1241]} = (x[1241]+y[1241]+z[1241]);
assign {c[1243],s[1242]} = (x[1242]+y[1242]+z[1242]);
assign {c[1244],s[1243]} = (x[1243]+y[1243]+z[1243]);
assign {c[1245],s[1244]} = (x[1244]+y[1244]+z[1244]);
assign {c[1246],s[1245]} = (x[1245]+y[1245]+z[1245]);
assign {c[1247],s[1246]} = (x[1246]+y[1246]+z[1246]);
assign {c[1248],s[1247]} = (x[1247]+y[1247]+z[1247]);
assign {c[1249],s[1248]} = (x[1248]+y[1248]+z[1248]);
assign {c[1250],s[1249]} = (x[1249]+y[1249]+z[1249]);
assign {c[1251],s[1250]} = (x[1250]+y[1250]+z[1250]);
assign {c[1252],s[1251]} = (x[1251]+y[1251]+z[1251]);
assign {c[1253],s[1252]} = (x[1252]+y[1252]+z[1252]);
assign {c[1254],s[1253]} = (x[1253]+y[1253]+z[1253]);
assign {c[1255],s[1254]} = (x[1254]+y[1254]+z[1254]);
assign {c[1256],s[1255]} = (x[1255]+y[1255]+z[1255]);
assign {c[1257],s[1256]} = (x[1256]+y[1256]+z[1256]);
assign {c[1258],s[1257]} = (x[1257]+y[1257]+z[1257]);
assign {c[1259],s[1258]} = (x[1258]+y[1258]+z[1258]);
assign {c[1260],s[1259]} = (x[1259]+y[1259]+z[1259]);
assign {c[1261],s[1260]} = (x[1260]+y[1260]+z[1260]);
assign {c[1262],s[1261]} = (x[1261]+y[1261]+z[1261]);
assign {c[1263],s[1262]} = (x[1262]+y[1262]+z[1262]);
assign {c[1264],s[1263]} = (x[1263]+y[1263]+z[1263]);
assign {c[1265],s[1264]} = (x[1264]+y[1264]+z[1264]);
assign {c[1266],s[1265]} = (x[1265]+y[1265]+z[1265]);
assign {c[1267],s[1266]} = (x[1266]+y[1266]+z[1266]);
assign {c[1268],s[1267]} = (x[1267]+y[1267]+z[1267]);
assign {c[1269],s[1268]} = (x[1268]+y[1268]+z[1268]);
assign {c[1270],s[1269]} = (x[1269]+y[1269]+z[1269]);
assign {c[1271],s[1270]} = (x[1270]+y[1270]+z[1270]);
assign {c[1272],s[1271]} = (x[1271]+y[1271]+z[1271]);
assign {c[1273],s[1272]} = (x[1272]+y[1272]+z[1272]);
assign {c[1274],s[1273]} = (x[1273]+y[1273]+z[1273]);
assign {c[1275],s[1274]} = (x[1274]+y[1274]+z[1274]);
assign {c[1276],s[1275]} = (x[1275]+y[1275]+z[1275]);
assign {c[1277],s[1276]} = (x[1276]+y[1276]+z[1276]);
assign {c[1278],s[1277]} = (x[1277]+y[1277]+z[1277]);
assign {c[1279],s[1278]} = (x[1278]+y[1278]+z[1278]);
assign {c[1280],s[1279]} = (x[1279]+y[1279]+z[1279]);
assign {c[1281],s[1280]} = (x[1280]+y[1280]+z[1280]);
assign {c[1282],s[1281]} = (x[1281]+y[1281]+z[1281]);
assign {c[1283],s[1282]} = (x[1282]+y[1282]+z[1282]);
assign {c[1284],s[1283]} = (x[1283]+y[1283]+z[1283]);
assign {c[1285],s[1284]} = (x[1284]+y[1284]+z[1284]);
assign {c[1286],s[1285]} = (x[1285]+y[1285]+z[1285]);
assign {c[1287],s[1286]} = (x[1286]+y[1286]+z[1286]);
assign {c[1288],s[1287]} = (x[1287]+y[1287]+z[1287]);
assign {c[1289],s[1288]} = (x[1288]+y[1288]+z[1288]);
assign {c[1290],s[1289]} = (x[1289]+y[1289]+z[1289]);
assign {c[1291],s[1290]} = (x[1290]+y[1290]+z[1290]);
assign {c[1292],s[1291]} = (x[1291]+y[1291]+z[1291]);
assign {c[1293],s[1292]} = (x[1292]+y[1292]+z[1292]);
assign {c[1294],s[1293]} = (x[1293]+y[1293]+z[1293]);
assign {c[1295],s[1294]} = (x[1294]+y[1294]+z[1294]);
assign {c[1296],s[1295]} = (x[1295]+y[1295]+z[1295]);
assign {c[1297],s[1296]} = (x[1296]+y[1296]+z[1296]);
assign {c[1298],s[1297]} = (x[1297]+y[1297]+z[1297]);
assign {c[1299],s[1298]} = (x[1298]+y[1298]+z[1298]);
assign {c[1300],s[1299]} = (x[1299]+y[1299]+z[1299]);
assign {c[1301],s[1300]} = (x[1300]+y[1300]+z[1300]);
assign {c[1302],s[1301]} = (x[1301]+y[1301]+z[1301]);
assign {c[1303],s[1302]} = (x[1302]+y[1302]+z[1302]);
assign {c[1304],s[1303]} = (x[1303]+y[1303]+z[1303]);
assign {c[1305],s[1304]} = (x[1304]+y[1304]+z[1304]);
assign {c[1306],s[1305]} = (x[1305]+y[1305]+z[1305]);
assign {c[1307],s[1306]} = (x[1306]+y[1306]+z[1306]);
assign {c[1308],s[1307]} = (x[1307]+y[1307]+z[1307]);
assign {c[1309],s[1308]} = (x[1308]+y[1308]+z[1308]);
assign {c[1310],s[1309]} = (x[1309]+y[1309]+z[1309]);
assign {c[1311],s[1310]} = (x[1310]+y[1310]+z[1310]);
assign {c[1312],s[1311]} = (x[1311]+y[1311]+z[1311]);
assign {c[1313],s[1312]} = (x[1312]+y[1312]+z[1312]);
assign {c[1314],s[1313]} = (x[1313]+y[1313]+z[1313]);
assign {c[1315],s[1314]} = (x[1314]+y[1314]+z[1314]);
assign {c[1316],s[1315]} = (x[1315]+y[1315]+z[1315]);
assign {c[1317],s[1316]} = (x[1316]+y[1316]+z[1316]);
assign {c[1318],s[1317]} = (x[1317]+y[1317]+z[1317]);
assign {c[1319],s[1318]} = (x[1318]+y[1318]+z[1318]);
assign {c[1320],s[1319]} = (x[1319]+y[1319]+z[1319]);
assign {c[1321],s[1320]} = (x[1320]+y[1320]+z[1320]);
assign {c[1322],s[1321]} = (x[1321]+y[1321]+z[1321]);
assign {c[1323],s[1322]} = (x[1322]+y[1322]+z[1322]);
assign {c[1324],s[1323]} = (x[1323]+y[1323]+z[1323]);
assign {c[1325],s[1324]} = (x[1324]+y[1324]+z[1324]);
assign {c[1326],s[1325]} = (x[1325]+y[1325]+z[1325]);
assign {c[1327],s[1326]} = (x[1326]+y[1326]+z[1326]);
assign {c[1328],s[1327]} = (x[1327]+y[1327]+z[1327]);
assign {c[1329],s[1328]} = (x[1328]+y[1328]+z[1328]);
assign {c[1330],s[1329]} = (x[1329]+y[1329]+z[1329]);
assign {c[1331],s[1330]} = (x[1330]+y[1330]+z[1330]);
assign {c[1332],s[1331]} = (x[1331]+y[1331]+z[1331]);
assign {c[1333],s[1332]} = (x[1332]+y[1332]+z[1332]);
assign {c[1334],s[1333]} = (x[1333]+y[1333]+z[1333]);
assign {c[1335],s[1334]} = (x[1334]+y[1334]+z[1334]);
assign {c[1336],s[1335]} = (x[1335]+y[1335]+z[1335]);
assign {c[1337],s[1336]} = (x[1336]+y[1336]+z[1336]);
assign {c[1338],s[1337]} = (x[1337]+y[1337]+z[1337]);
assign {c[1339],s[1338]} = (x[1338]+y[1338]+z[1338]);
assign {c[1340],s[1339]} = (x[1339]+y[1339]+z[1339]);
assign {c[1341],s[1340]} = (x[1340]+y[1340]+z[1340]);
assign {c[1342],s[1341]} = (x[1341]+y[1341]+z[1341]);
assign {c[1343],s[1342]} = (x[1342]+y[1342]+z[1342]);
assign {c[1344],s[1343]} = (x[1343]+y[1343]+z[1343]);
assign {c[1345],s[1344]} = (x[1344]+y[1344]+z[1344]);
assign {c[1346],s[1345]} = (x[1345]+y[1345]+z[1345]);
assign {c[1347],s[1346]} = (x[1346]+y[1346]+z[1346]);
assign {c[1348],s[1347]} = (x[1347]+y[1347]+z[1347]);
assign {c[1349],s[1348]} = (x[1348]+y[1348]+z[1348]);
assign {c[1350],s[1349]} = (x[1349]+y[1349]+z[1349]);
assign {c[1351],s[1350]} = (x[1350]+y[1350]+z[1350]);
assign {c[1352],s[1351]} = (x[1351]+y[1351]+z[1351]);
assign {c[1353],s[1352]} = (x[1352]+y[1352]+z[1352]);
assign {c[1354],s[1353]} = (x[1353]+y[1353]+z[1353]);
assign {c[1355],s[1354]} = (x[1354]+y[1354]+z[1354]);
assign {c[1356],s[1355]} = (x[1355]+y[1355]+z[1355]);
assign {c[1357],s[1356]} = (x[1356]+y[1356]+z[1356]);
assign {c[1358],s[1357]} = (x[1357]+y[1357]+z[1357]);
assign {c[1359],s[1358]} = (x[1358]+y[1358]+z[1358]);
assign {c[1360],s[1359]} = (x[1359]+y[1359]+z[1359]);
assign {c[1361],s[1360]} = (x[1360]+y[1360]+z[1360]);
assign {c[1362],s[1361]} = (x[1361]+y[1361]+z[1361]);
assign {c[1363],s[1362]} = (x[1362]+y[1362]+z[1362]);
assign {c[1364],s[1363]} = (x[1363]+y[1363]+z[1363]);
assign {c[1365],s[1364]} = (x[1364]+y[1364]+z[1364]);
assign {c[1366],s[1365]} = (x[1365]+y[1365]+z[1365]);
assign {c[1367],s[1366]} = (x[1366]+y[1366]+z[1366]);
assign {c[1368],s[1367]} = (x[1367]+y[1367]+z[1367]);
assign {c[1369],s[1368]} = (x[1368]+y[1368]+z[1368]);
assign {c[1370],s[1369]} = (x[1369]+y[1369]+z[1369]);
assign {c[1371],s[1370]} = (x[1370]+y[1370]+z[1370]);
assign {c[1372],s[1371]} = (x[1371]+y[1371]+z[1371]);
assign {c[1373],s[1372]} = (x[1372]+y[1372]+z[1372]);
assign {c[1374],s[1373]} = (x[1373]+y[1373]+z[1373]);
assign {c[1375],s[1374]} = (x[1374]+y[1374]+z[1374]);
assign {c[1376],s[1375]} = (x[1375]+y[1375]+z[1375]);
assign {c[1377],s[1376]} = (x[1376]+y[1376]+z[1376]);
assign {c[1378],s[1377]} = (x[1377]+y[1377]+z[1377]);
assign {c[1379],s[1378]} = (x[1378]+y[1378]+z[1378]);
assign {c[1380],s[1379]} = (x[1379]+y[1379]+z[1379]);
assign {c[1381],s[1380]} = (x[1380]+y[1380]+z[1380]);
assign {c[1382],s[1381]} = (x[1381]+y[1381]+z[1381]);
assign {c[1383],s[1382]} = (x[1382]+y[1382]+z[1382]);
assign {c[1384],s[1383]} = (x[1383]+y[1383]+z[1383]);
assign {c[1385],s[1384]} = (x[1384]+y[1384]+z[1384]);
assign {c[1386],s[1385]} = (x[1385]+y[1385]+z[1385]);
assign {c[1387],s[1386]} = (x[1386]+y[1386]+z[1386]);
assign {c[1388],s[1387]} = (x[1387]+y[1387]+z[1387]);
assign {c[1389],s[1388]} = (x[1388]+y[1388]+z[1388]);
assign {c[1390],s[1389]} = (x[1389]+y[1389]+z[1389]);
assign {c[1391],s[1390]} = (x[1390]+y[1390]+z[1390]);
assign {c[1392],s[1391]} = (x[1391]+y[1391]+z[1391]);
assign {c[1393],s[1392]} = (x[1392]+y[1392]+z[1392]);
assign {c[1394],s[1393]} = (x[1393]+y[1393]+z[1393]);
assign {c[1395],s[1394]} = (x[1394]+y[1394]+z[1394]);
assign {c[1396],s[1395]} = (x[1395]+y[1395]+z[1395]);
assign {c[1397],s[1396]} = (x[1396]+y[1396]+z[1396]);
assign {c[1398],s[1397]} = (x[1397]+y[1397]+z[1397]);
assign {c[1399],s[1398]} = (x[1398]+y[1398]+z[1398]);
assign {c[1400],s[1399]} = (x[1399]+y[1399]+z[1399]);
assign {c[1401],s[1400]} = (x[1400]+y[1400]+z[1400]);
assign {c[1402],s[1401]} = (x[1401]+y[1401]+z[1401]);
assign {c[1403],s[1402]} = (x[1402]+y[1402]+z[1402]);
assign {c[1404],s[1403]} = (x[1403]+y[1403]+z[1403]);
assign {c[1405],s[1404]} = (x[1404]+y[1404]+z[1404]);
assign {c[1406],s[1405]} = (x[1405]+y[1405]+z[1405]);
assign {c[1407],s[1406]} = (x[1406]+y[1406]+z[1406]);
assign {c[1408],s[1407]} = (x[1407]+y[1407]+z[1407]);
assign {c[1409],s[1408]} = (x[1408]+y[1408]+z[1408]);
assign {c[1410],s[1409]} = (x[1409]+y[1409]+z[1409]);
assign {c[1411],s[1410]} = (x[1410]+y[1410]+z[1410]);
assign {c[1412],s[1411]} = (x[1411]+y[1411]+z[1411]);
assign {c[1413],s[1412]} = (x[1412]+y[1412]+z[1412]);
assign {c[1414],s[1413]} = (x[1413]+y[1413]+z[1413]);
assign {c[1415],s[1414]} = (x[1414]+y[1414]+z[1414]);
assign {c[1416],s[1415]} = (x[1415]+y[1415]+z[1415]);
assign {c[1417],s[1416]} = (x[1416]+y[1416]+z[1416]);
assign {c[1418],s[1417]} = (x[1417]+y[1417]+z[1417]);
assign {c[1419],s[1418]} = (x[1418]+y[1418]+z[1418]);
assign {c[1420],s[1419]} = (x[1419]+y[1419]+z[1419]);
assign {c[1421],s[1420]} = (x[1420]+y[1420]+z[1420]);
assign {c[1422],s[1421]} = (x[1421]+y[1421]+z[1421]);
assign {c[1423],s[1422]} = (x[1422]+y[1422]+z[1422]);
assign {c[1424],s[1423]} = (x[1423]+y[1423]+z[1423]);
assign {c[1425],s[1424]} = (x[1424]+y[1424]+z[1424]);
assign {c[1426],s[1425]} = (x[1425]+y[1425]+z[1425]);
assign {c[1427],s[1426]} = (x[1426]+y[1426]+z[1426]);
assign {c[1428],s[1427]} = (x[1427]+y[1427]+z[1427]);
assign {c[1429],s[1428]} = (x[1428]+y[1428]+z[1428]);
assign {c[1430],s[1429]} = (x[1429]+y[1429]+z[1429]);
assign {c[1431],s[1430]} = (x[1430]+y[1430]+z[1430]);
assign {c[1432],s[1431]} = (x[1431]+y[1431]+z[1431]);
assign {c[1433],s[1432]} = (x[1432]+y[1432]+z[1432]);
assign {c[1434],s[1433]} = (x[1433]+y[1433]+z[1433]);
assign {c[1435],s[1434]} = (x[1434]+y[1434]+z[1434]);
assign {c[1436],s[1435]} = (x[1435]+y[1435]+z[1435]);
assign {c[1437],s[1436]} = (x[1436]+y[1436]+z[1436]);
assign {c[1438],s[1437]} = (x[1437]+y[1437]+z[1437]);
assign {c[1439],s[1438]} = (x[1438]+y[1438]+z[1438]);
assign {c[1440],s[1439]} = (x[1439]+y[1439]+z[1439]);
assign {c[1441],s[1440]} = (x[1440]+y[1440]+z[1440]);
assign {c[1442],s[1441]} = (x[1441]+y[1441]+z[1441]);
assign {c[1443],s[1442]} = (x[1442]+y[1442]+z[1442]);
assign {c[1444],s[1443]} = (x[1443]+y[1443]+z[1443]);
assign {c[1445],s[1444]} = (x[1444]+y[1444]+z[1444]);
assign {c[1446],s[1445]} = (x[1445]+y[1445]+z[1445]);
assign {c[1447],s[1446]} = (x[1446]+y[1446]+z[1446]);
assign {c[1448],s[1447]} = (x[1447]+y[1447]+z[1447]);
assign {c[1449],s[1448]} = (x[1448]+y[1448]+z[1448]);
assign {c[1450],s[1449]} = (x[1449]+y[1449]+z[1449]);
assign {c[1451],s[1450]} = (x[1450]+y[1450]+z[1450]);
assign {c[1452],s[1451]} = (x[1451]+y[1451]+z[1451]);
assign {c[1453],s[1452]} = (x[1452]+y[1452]+z[1452]);
assign {c[1454],s[1453]} = (x[1453]+y[1453]+z[1453]);
assign {c[1455],s[1454]} = (x[1454]+y[1454]+z[1454]);
assign {c[1456],s[1455]} = (x[1455]+y[1455]+z[1455]);
assign {c[1457],s[1456]} = (x[1456]+y[1456]+z[1456]);
assign {c[1458],s[1457]} = (x[1457]+y[1457]+z[1457]);
assign {c[1459],s[1458]} = (x[1458]+y[1458]+z[1458]);
assign {c[1460],s[1459]} = (x[1459]+y[1459]+z[1459]);
assign {c[1461],s[1460]} = (x[1460]+y[1460]+z[1460]);
assign {c[1462],s[1461]} = (x[1461]+y[1461]+z[1461]);
assign {c[1463],s[1462]} = (x[1462]+y[1462]+z[1462]);
assign {c[1464],s[1463]} = (x[1463]+y[1463]+z[1463]);
assign {c[1465],s[1464]} = (x[1464]+y[1464]+z[1464]);
assign {c[1466],s[1465]} = (x[1465]+y[1465]+z[1465]);
assign {c[1467],s[1466]} = (x[1466]+y[1466]+z[1466]);
assign {c[1468],s[1467]} = (x[1467]+y[1467]+z[1467]);
assign {c[1469],s[1468]} = (x[1468]+y[1468]+z[1468]);
assign {c[1470],s[1469]} = (x[1469]+y[1469]+z[1469]);
assign {c[1471],s[1470]} = (x[1470]+y[1470]+z[1470]);
assign {c[1472],s[1471]} = (x[1471]+y[1471]+z[1471]);
assign {c[1473],s[1472]} = (x[1472]+y[1472]+z[1472]);
assign {c[1474],s[1473]} = (x[1473]+y[1473]+z[1473]);
assign {c[1475],s[1474]} = (x[1474]+y[1474]+z[1474]);
assign {c[1476],s[1475]} = (x[1475]+y[1475]+z[1475]);
assign {c[1477],s[1476]} = (x[1476]+y[1476]+z[1476]);
assign {c[1478],s[1477]} = (x[1477]+y[1477]+z[1477]);
assign {c[1479],s[1478]} = (x[1478]+y[1478]+z[1478]);
assign {c[1480],s[1479]} = (x[1479]+y[1479]+z[1479]);
assign {c[1481],s[1480]} = (x[1480]+y[1480]+z[1480]);
assign {c[1482],s[1481]} = (x[1481]+y[1481]+z[1481]);
assign {c[1483],s[1482]} = (x[1482]+y[1482]+z[1482]);
assign {c[1484],s[1483]} = (x[1483]+y[1483]+z[1483]);
assign {c[1485],s[1484]} = (x[1484]+y[1484]+z[1484]);
assign {c[1486],s[1485]} = (x[1485]+y[1485]+z[1485]);
assign {c[1487],s[1486]} = (x[1486]+y[1486]+z[1486]);
assign {c[1488],s[1487]} = (x[1487]+y[1487]+z[1487]);
assign {c[1489],s[1488]} = (x[1488]+y[1488]+z[1488]);
assign {c[1490],s[1489]} = (x[1489]+y[1489]+z[1489]);
assign {c[1491],s[1490]} = (x[1490]+y[1490]+z[1490]);
assign {c[1492],s[1491]} = (x[1491]+y[1491]+z[1491]);
assign {c[1493],s[1492]} = (x[1492]+y[1492]+z[1492]);
assign {c[1494],s[1493]} = (x[1493]+y[1493]+z[1493]);
assign {c[1495],s[1494]} = (x[1494]+y[1494]+z[1494]);
assign {c[1496],s[1495]} = (x[1495]+y[1495]+z[1495]);
assign {c[1497],s[1496]} = (x[1496]+y[1496]+z[1496]);
assign {c[1498],s[1497]} = (x[1497]+y[1497]+z[1497]);
assign {c[1499],s[1498]} = (x[1498]+y[1498]+z[1498]);
assign {c[1500],s[1499]} = (x[1499]+y[1499]+z[1499]);
assign {c[1501],s[1500]} = (x[1500]+y[1500]+z[1500]);
assign {c[1502],s[1501]} = (x[1501]+y[1501]+z[1501]);
assign {c[1503],s[1502]} = (x[1502]+y[1502]+z[1502]);
assign {c[1504],s[1503]} = (x[1503]+y[1503]+z[1503]);
assign {c[1505],s[1504]} = (x[1504]+y[1504]+z[1504]);
assign {c[1506],s[1505]} = (x[1505]+y[1505]+z[1505]);
assign {c[1507],s[1506]} = (x[1506]+y[1506]+z[1506]);
assign {c[1508],s[1507]} = (x[1507]+y[1507]+z[1507]);
assign {c[1509],s[1508]} = (x[1508]+y[1508]+z[1508]);
assign {dummy,s[1509]} = (x[1509]+y[1509]+z[1509]);

endmodule
    