

module csa_tree_1509x1509_truncated(
    input [2277080:0] A, // lines are appended together
    output[1508:0] B_0,
    output[1508:0] B_1
);

wire [1518053:0] tree_1;
wire [1012538:0] tree_2;
wire [676031:0] tree_3;
wire [451190:0] tree_4;
wire [301799:0] tree_5;
wire [202205:0] tree_6;
wire [135809:0] tree_7;
wire [90539:0] tree_8;
wire [60359:0] tree_9;
wire [40742:0] tree_10;
wire [27161:0] tree_11;
wire [18107:0] tree_12;
wire [12071:0] tree_13;
wire [9053:0] tree_14;
wire [6035:0] tree_15;
wire [4526:0] tree_16;
wire [3017:0] tree_17;
// layer-1
csa_1509 csau_1509_i0(A[1508:0],A[3017:1509],A[4526:3018],tree_1[1508:0],tree_1[3017:1509]);
csa_1509 csau_1509_i1(A[6035:4527],A[7544:6036],A[9053:7545],tree_1[4526:3018],tree_1[6035:4527]);
csa_1509 csau_1509_i2(A[10562:9054],A[12071:10563],A[13580:12072],tree_1[7544:6036],tree_1[9053:7545]);
csa_1509 csau_1509_i3(A[15089:13581],A[16598:15090],A[18107:16599],tree_1[10562:9054],tree_1[12071:10563]);
csa_1509 csau_1509_i4(A[19616:18108],A[21125:19617],A[22634:21126],tree_1[13580:12072],tree_1[15089:13581]);
csa_1509 csau_1509_i5(A[24143:22635],A[25652:24144],A[27161:25653],tree_1[16598:15090],tree_1[18107:16599]);
csa_1509 csau_1509_i6(A[28670:27162],A[30179:28671],A[31688:30180],tree_1[19616:18108],tree_1[21125:19617]);
csa_1509 csau_1509_i7(A[33197:31689],A[34706:33198],A[36215:34707],tree_1[22634:21126],tree_1[24143:22635]);
csa_1509 csau_1509_i8(A[37724:36216],A[39233:37725],A[40742:39234],tree_1[25652:24144],tree_1[27161:25653]);
csa_1509 csau_1509_i9(A[42251:40743],A[43760:42252],A[45269:43761],tree_1[28670:27162],tree_1[30179:28671]);
csa_1509 csau_1509_i10(A[46778:45270],A[48287:46779],A[49796:48288],tree_1[31688:30180],tree_1[33197:31689]);
csa_1509 csau_1509_i11(A[51305:49797],A[52814:51306],A[54323:52815],tree_1[34706:33198],tree_1[36215:34707]);
csa_1509 csau_1509_i12(A[55832:54324],A[57341:55833],A[58850:57342],tree_1[37724:36216],tree_1[39233:37725]);
csa_1509 csau_1509_i13(A[60359:58851],A[61868:60360],A[63377:61869],tree_1[40742:39234],tree_1[42251:40743]);
csa_1509 csau_1509_i14(A[64886:63378],A[66395:64887],A[67904:66396],tree_1[43760:42252],tree_1[45269:43761]);
csa_1509 csau_1509_i15(A[69413:67905],A[70922:69414],A[72431:70923],tree_1[46778:45270],tree_1[48287:46779]);
csa_1509 csau_1509_i16(A[73940:72432],A[75449:73941],A[76958:75450],tree_1[49796:48288],tree_1[51305:49797]);
csa_1509 csau_1509_i17(A[78467:76959],A[79976:78468],A[81485:79977],tree_1[52814:51306],tree_1[54323:52815]);
csa_1509 csau_1509_i18(A[82994:81486],A[84503:82995],A[86012:84504],tree_1[55832:54324],tree_1[57341:55833]);
csa_1509 csau_1509_i19(A[87521:86013],A[89030:87522],A[90539:89031],tree_1[58850:57342],tree_1[60359:58851]);
csa_1509 csau_1509_i20(A[92048:90540],A[93557:92049],A[95066:93558],tree_1[61868:60360],tree_1[63377:61869]);
csa_1509 csau_1509_i21(A[96575:95067],A[98084:96576],A[99593:98085],tree_1[64886:63378],tree_1[66395:64887]);
csa_1509 csau_1509_i22(A[101102:99594],A[102611:101103],A[104120:102612],tree_1[67904:66396],tree_1[69413:67905]);
csa_1509 csau_1509_i23(A[105629:104121],A[107138:105630],A[108647:107139],tree_1[70922:69414],tree_1[72431:70923]);
csa_1509 csau_1509_i24(A[110156:108648],A[111665:110157],A[113174:111666],tree_1[73940:72432],tree_1[75449:73941]);
csa_1509 csau_1509_i25(A[114683:113175],A[116192:114684],A[117701:116193],tree_1[76958:75450],tree_1[78467:76959]);
csa_1509 csau_1509_i26(A[119210:117702],A[120719:119211],A[122228:120720],tree_1[79976:78468],tree_1[81485:79977]);
csa_1509 csau_1509_i27(A[123737:122229],A[125246:123738],A[126755:125247],tree_1[82994:81486],tree_1[84503:82995]);
csa_1509 csau_1509_i28(A[128264:126756],A[129773:128265],A[131282:129774],tree_1[86012:84504],tree_1[87521:86013]);
csa_1509 csau_1509_i29(A[132791:131283],A[134300:132792],A[135809:134301],tree_1[89030:87522],tree_1[90539:89031]);
csa_1509 csau_1509_i30(A[137318:135810],A[138827:137319],A[140336:138828],tree_1[92048:90540],tree_1[93557:92049]);
csa_1509 csau_1509_i31(A[141845:140337],A[143354:141846],A[144863:143355],tree_1[95066:93558],tree_1[96575:95067]);
csa_1509 csau_1509_i32(A[146372:144864],A[147881:146373],A[149390:147882],tree_1[98084:96576],tree_1[99593:98085]);
csa_1509 csau_1509_i33(A[150899:149391],A[152408:150900],A[153917:152409],tree_1[101102:99594],tree_1[102611:101103]);
csa_1509 csau_1509_i34(A[155426:153918],A[156935:155427],A[158444:156936],tree_1[104120:102612],tree_1[105629:104121]);
csa_1509 csau_1509_i35(A[159953:158445],A[161462:159954],A[162971:161463],tree_1[107138:105630],tree_1[108647:107139]);
csa_1509 csau_1509_i36(A[164480:162972],A[165989:164481],A[167498:165990],tree_1[110156:108648],tree_1[111665:110157]);
csa_1509 csau_1509_i37(A[169007:167499],A[170516:169008],A[172025:170517],tree_1[113174:111666],tree_1[114683:113175]);
csa_1509 csau_1509_i38(A[173534:172026],A[175043:173535],A[176552:175044],tree_1[116192:114684],tree_1[117701:116193]);
csa_1509 csau_1509_i39(A[178061:176553],A[179570:178062],A[181079:179571],tree_1[119210:117702],tree_1[120719:119211]);
csa_1509 csau_1509_i40(A[182588:181080],A[184097:182589],A[185606:184098],tree_1[122228:120720],tree_1[123737:122229]);
csa_1509 csau_1509_i41(A[187115:185607],A[188624:187116],A[190133:188625],tree_1[125246:123738],tree_1[126755:125247]);
csa_1509 csau_1509_i42(A[191642:190134],A[193151:191643],A[194660:193152],tree_1[128264:126756],tree_1[129773:128265]);
csa_1509 csau_1509_i43(A[196169:194661],A[197678:196170],A[199187:197679],tree_1[131282:129774],tree_1[132791:131283]);
csa_1509 csau_1509_i44(A[200696:199188],A[202205:200697],A[203714:202206],tree_1[134300:132792],tree_1[135809:134301]);
csa_1509 csau_1509_i45(A[205223:203715],A[206732:205224],A[208241:206733],tree_1[137318:135810],tree_1[138827:137319]);
csa_1509 csau_1509_i46(A[209750:208242],A[211259:209751],A[212768:211260],tree_1[140336:138828],tree_1[141845:140337]);
csa_1509 csau_1509_i47(A[214277:212769],A[215786:214278],A[217295:215787],tree_1[143354:141846],tree_1[144863:143355]);
csa_1509 csau_1509_i48(A[218804:217296],A[220313:218805],A[221822:220314],tree_1[146372:144864],tree_1[147881:146373]);
csa_1509 csau_1509_i49(A[223331:221823],A[224840:223332],A[226349:224841],tree_1[149390:147882],tree_1[150899:149391]);
csa_1509 csau_1509_i50(A[227858:226350],A[229367:227859],A[230876:229368],tree_1[152408:150900],tree_1[153917:152409]);
csa_1509 csau_1509_i51(A[232385:230877],A[233894:232386],A[235403:233895],tree_1[155426:153918],tree_1[156935:155427]);
csa_1509 csau_1509_i52(A[236912:235404],A[238421:236913],A[239930:238422],tree_1[158444:156936],tree_1[159953:158445]);
csa_1509 csau_1509_i53(A[241439:239931],A[242948:241440],A[244457:242949],tree_1[161462:159954],tree_1[162971:161463]);
csa_1509 csau_1509_i54(A[245966:244458],A[247475:245967],A[248984:247476],tree_1[164480:162972],tree_1[165989:164481]);
csa_1509 csau_1509_i55(A[250493:248985],A[252002:250494],A[253511:252003],tree_1[167498:165990],tree_1[169007:167499]);
csa_1509 csau_1509_i56(A[255020:253512],A[256529:255021],A[258038:256530],tree_1[170516:169008],tree_1[172025:170517]);
csa_1509 csau_1509_i57(A[259547:258039],A[261056:259548],A[262565:261057],tree_1[173534:172026],tree_1[175043:173535]);
csa_1509 csau_1509_i58(A[264074:262566],A[265583:264075],A[267092:265584],tree_1[176552:175044],tree_1[178061:176553]);
csa_1509 csau_1509_i59(A[268601:267093],A[270110:268602],A[271619:270111],tree_1[179570:178062],tree_1[181079:179571]);
csa_1509 csau_1509_i60(A[273128:271620],A[274637:273129],A[276146:274638],tree_1[182588:181080],tree_1[184097:182589]);
csa_1509 csau_1509_i61(A[277655:276147],A[279164:277656],A[280673:279165],tree_1[185606:184098],tree_1[187115:185607]);
csa_1509 csau_1509_i62(A[282182:280674],A[283691:282183],A[285200:283692],tree_1[188624:187116],tree_1[190133:188625]);
csa_1509 csau_1509_i63(A[286709:285201],A[288218:286710],A[289727:288219],tree_1[191642:190134],tree_1[193151:191643]);
csa_1509 csau_1509_i64(A[291236:289728],A[292745:291237],A[294254:292746],tree_1[194660:193152],tree_1[196169:194661]);
csa_1509 csau_1509_i65(A[295763:294255],A[297272:295764],A[298781:297273],tree_1[197678:196170],tree_1[199187:197679]);
csa_1509 csau_1509_i66(A[300290:298782],A[301799:300291],A[303308:301800],tree_1[200696:199188],tree_1[202205:200697]);
csa_1509 csau_1509_i67(A[304817:303309],A[306326:304818],A[307835:306327],tree_1[203714:202206],tree_1[205223:203715]);
csa_1509 csau_1509_i68(A[309344:307836],A[310853:309345],A[312362:310854],tree_1[206732:205224],tree_1[208241:206733]);
csa_1509 csau_1509_i69(A[313871:312363],A[315380:313872],A[316889:315381],tree_1[209750:208242],tree_1[211259:209751]);
csa_1509 csau_1509_i70(A[318398:316890],A[319907:318399],A[321416:319908],tree_1[212768:211260],tree_1[214277:212769]);
csa_1509 csau_1509_i71(A[322925:321417],A[324434:322926],A[325943:324435],tree_1[215786:214278],tree_1[217295:215787]);
csa_1509 csau_1509_i72(A[327452:325944],A[328961:327453],A[330470:328962],tree_1[218804:217296],tree_1[220313:218805]);
csa_1509 csau_1509_i73(A[331979:330471],A[333488:331980],A[334997:333489],tree_1[221822:220314],tree_1[223331:221823]);
csa_1509 csau_1509_i74(A[336506:334998],A[338015:336507],A[339524:338016],tree_1[224840:223332],tree_1[226349:224841]);
csa_1509 csau_1509_i75(A[341033:339525],A[342542:341034],A[344051:342543],tree_1[227858:226350],tree_1[229367:227859]);
csa_1509 csau_1509_i76(A[345560:344052],A[347069:345561],A[348578:347070],tree_1[230876:229368],tree_1[232385:230877]);
csa_1509 csau_1509_i77(A[350087:348579],A[351596:350088],A[353105:351597],tree_1[233894:232386],tree_1[235403:233895]);
csa_1509 csau_1509_i78(A[354614:353106],A[356123:354615],A[357632:356124],tree_1[236912:235404],tree_1[238421:236913]);
csa_1509 csau_1509_i79(A[359141:357633],A[360650:359142],A[362159:360651],tree_1[239930:238422],tree_1[241439:239931]);
csa_1509 csau_1509_i80(A[363668:362160],A[365177:363669],A[366686:365178],tree_1[242948:241440],tree_1[244457:242949]);
csa_1509 csau_1509_i81(A[368195:366687],A[369704:368196],A[371213:369705],tree_1[245966:244458],tree_1[247475:245967]);
csa_1509 csau_1509_i82(A[372722:371214],A[374231:372723],A[375740:374232],tree_1[248984:247476],tree_1[250493:248985]);
csa_1509 csau_1509_i83(A[377249:375741],A[378758:377250],A[380267:378759],tree_1[252002:250494],tree_1[253511:252003]);
csa_1509 csau_1509_i84(A[381776:380268],A[383285:381777],A[384794:383286],tree_1[255020:253512],tree_1[256529:255021]);
csa_1509 csau_1509_i85(A[386303:384795],A[387812:386304],A[389321:387813],tree_1[258038:256530],tree_1[259547:258039]);
csa_1509 csau_1509_i86(A[390830:389322],A[392339:390831],A[393848:392340],tree_1[261056:259548],tree_1[262565:261057]);
csa_1509 csau_1509_i87(A[395357:393849],A[396866:395358],A[398375:396867],tree_1[264074:262566],tree_1[265583:264075]);
csa_1509 csau_1509_i88(A[399884:398376],A[401393:399885],A[402902:401394],tree_1[267092:265584],tree_1[268601:267093]);
csa_1509 csau_1509_i89(A[404411:402903],A[405920:404412],A[407429:405921],tree_1[270110:268602],tree_1[271619:270111]);
csa_1509 csau_1509_i90(A[408938:407430],A[410447:408939],A[411956:410448],tree_1[273128:271620],tree_1[274637:273129]);
csa_1509 csau_1509_i91(A[413465:411957],A[414974:413466],A[416483:414975],tree_1[276146:274638],tree_1[277655:276147]);
csa_1509 csau_1509_i92(A[417992:416484],A[419501:417993],A[421010:419502],tree_1[279164:277656],tree_1[280673:279165]);
csa_1509 csau_1509_i93(A[422519:421011],A[424028:422520],A[425537:424029],tree_1[282182:280674],tree_1[283691:282183]);
csa_1509 csau_1509_i94(A[427046:425538],A[428555:427047],A[430064:428556],tree_1[285200:283692],tree_1[286709:285201]);
csa_1509 csau_1509_i95(A[431573:430065],A[433082:431574],A[434591:433083],tree_1[288218:286710],tree_1[289727:288219]);
csa_1509 csau_1509_i96(A[436100:434592],A[437609:436101],A[439118:437610],tree_1[291236:289728],tree_1[292745:291237]);
csa_1509 csau_1509_i97(A[440627:439119],A[442136:440628],A[443645:442137],tree_1[294254:292746],tree_1[295763:294255]);
csa_1509 csau_1509_i98(A[445154:443646],A[446663:445155],A[448172:446664],tree_1[297272:295764],tree_1[298781:297273]);
csa_1509 csau_1509_i99(A[449681:448173],A[451190:449682],A[452699:451191],tree_1[300290:298782],tree_1[301799:300291]);
csa_1509 csau_1509_i100(A[454208:452700],A[455717:454209],A[457226:455718],tree_1[303308:301800],tree_1[304817:303309]);
csa_1509 csau_1509_i101(A[458735:457227],A[460244:458736],A[461753:460245],tree_1[306326:304818],tree_1[307835:306327]);
csa_1509 csau_1509_i102(A[463262:461754],A[464771:463263],A[466280:464772],tree_1[309344:307836],tree_1[310853:309345]);
csa_1509 csau_1509_i103(A[467789:466281],A[469298:467790],A[470807:469299],tree_1[312362:310854],tree_1[313871:312363]);
csa_1509 csau_1509_i104(A[472316:470808],A[473825:472317],A[475334:473826],tree_1[315380:313872],tree_1[316889:315381]);
csa_1509 csau_1509_i105(A[476843:475335],A[478352:476844],A[479861:478353],tree_1[318398:316890],tree_1[319907:318399]);
csa_1509 csau_1509_i106(A[481370:479862],A[482879:481371],A[484388:482880],tree_1[321416:319908],tree_1[322925:321417]);
csa_1509 csau_1509_i107(A[485897:484389],A[487406:485898],A[488915:487407],tree_1[324434:322926],tree_1[325943:324435]);
csa_1509 csau_1509_i108(A[490424:488916],A[491933:490425],A[493442:491934],tree_1[327452:325944],tree_1[328961:327453]);
csa_1509 csau_1509_i109(A[494951:493443],A[496460:494952],A[497969:496461],tree_1[330470:328962],tree_1[331979:330471]);
csa_1509 csau_1509_i110(A[499478:497970],A[500987:499479],A[502496:500988],tree_1[333488:331980],tree_1[334997:333489]);
csa_1509 csau_1509_i111(A[504005:502497],A[505514:504006],A[507023:505515],tree_1[336506:334998],tree_1[338015:336507]);
csa_1509 csau_1509_i112(A[508532:507024],A[510041:508533],A[511550:510042],tree_1[339524:338016],tree_1[341033:339525]);
csa_1509 csau_1509_i113(A[513059:511551],A[514568:513060],A[516077:514569],tree_1[342542:341034],tree_1[344051:342543]);
csa_1509 csau_1509_i114(A[517586:516078],A[519095:517587],A[520604:519096],tree_1[345560:344052],tree_1[347069:345561]);
csa_1509 csau_1509_i115(A[522113:520605],A[523622:522114],A[525131:523623],tree_1[348578:347070],tree_1[350087:348579]);
csa_1509 csau_1509_i116(A[526640:525132],A[528149:526641],A[529658:528150],tree_1[351596:350088],tree_1[353105:351597]);
csa_1509 csau_1509_i117(A[531167:529659],A[532676:531168],A[534185:532677],tree_1[354614:353106],tree_1[356123:354615]);
csa_1509 csau_1509_i118(A[535694:534186],A[537203:535695],A[538712:537204],tree_1[357632:356124],tree_1[359141:357633]);
csa_1509 csau_1509_i119(A[540221:538713],A[541730:540222],A[543239:541731],tree_1[360650:359142],tree_1[362159:360651]);
csa_1509 csau_1509_i120(A[544748:543240],A[546257:544749],A[547766:546258],tree_1[363668:362160],tree_1[365177:363669]);
csa_1509 csau_1509_i121(A[549275:547767],A[550784:549276],A[552293:550785],tree_1[366686:365178],tree_1[368195:366687]);
csa_1509 csau_1509_i122(A[553802:552294],A[555311:553803],A[556820:555312],tree_1[369704:368196],tree_1[371213:369705]);
csa_1509 csau_1509_i123(A[558329:556821],A[559838:558330],A[561347:559839],tree_1[372722:371214],tree_1[374231:372723]);
csa_1509 csau_1509_i124(A[562856:561348],A[564365:562857],A[565874:564366],tree_1[375740:374232],tree_1[377249:375741]);
csa_1509 csau_1509_i125(A[567383:565875],A[568892:567384],A[570401:568893],tree_1[378758:377250],tree_1[380267:378759]);
csa_1509 csau_1509_i126(A[571910:570402],A[573419:571911],A[574928:573420],tree_1[381776:380268],tree_1[383285:381777]);
csa_1509 csau_1509_i127(A[576437:574929],A[577946:576438],A[579455:577947],tree_1[384794:383286],tree_1[386303:384795]);
csa_1509 csau_1509_i128(A[580964:579456],A[582473:580965],A[583982:582474],tree_1[387812:386304],tree_1[389321:387813]);
csa_1509 csau_1509_i129(A[585491:583983],A[587000:585492],A[588509:587001],tree_1[390830:389322],tree_1[392339:390831]);
csa_1509 csau_1509_i130(A[590018:588510],A[591527:590019],A[593036:591528],tree_1[393848:392340],tree_1[395357:393849]);
csa_1509 csau_1509_i131(A[594545:593037],A[596054:594546],A[597563:596055],tree_1[396866:395358],tree_1[398375:396867]);
csa_1509 csau_1509_i132(A[599072:597564],A[600581:599073],A[602090:600582],tree_1[399884:398376],tree_1[401393:399885]);
csa_1509 csau_1509_i133(A[603599:602091],A[605108:603600],A[606617:605109],tree_1[402902:401394],tree_1[404411:402903]);
csa_1509 csau_1509_i134(A[608126:606618],A[609635:608127],A[611144:609636],tree_1[405920:404412],tree_1[407429:405921]);
csa_1509 csau_1509_i135(A[612653:611145],A[614162:612654],A[615671:614163],tree_1[408938:407430],tree_1[410447:408939]);
csa_1509 csau_1509_i136(A[617180:615672],A[618689:617181],A[620198:618690],tree_1[411956:410448],tree_1[413465:411957]);
csa_1509 csau_1509_i137(A[621707:620199],A[623216:621708],A[624725:623217],tree_1[414974:413466],tree_1[416483:414975]);
csa_1509 csau_1509_i138(A[626234:624726],A[627743:626235],A[629252:627744],tree_1[417992:416484],tree_1[419501:417993]);
csa_1509 csau_1509_i139(A[630761:629253],A[632270:630762],A[633779:632271],tree_1[421010:419502],tree_1[422519:421011]);
csa_1509 csau_1509_i140(A[635288:633780],A[636797:635289],A[638306:636798],tree_1[424028:422520],tree_1[425537:424029]);
csa_1509 csau_1509_i141(A[639815:638307],A[641324:639816],A[642833:641325],tree_1[427046:425538],tree_1[428555:427047]);
csa_1509 csau_1509_i142(A[644342:642834],A[645851:644343],A[647360:645852],tree_1[430064:428556],tree_1[431573:430065]);
csa_1509 csau_1509_i143(A[648869:647361],A[650378:648870],A[651887:650379],tree_1[433082:431574],tree_1[434591:433083]);
csa_1509 csau_1509_i144(A[653396:651888],A[654905:653397],A[656414:654906],tree_1[436100:434592],tree_1[437609:436101]);
csa_1509 csau_1509_i145(A[657923:656415],A[659432:657924],A[660941:659433],tree_1[439118:437610],tree_1[440627:439119]);
csa_1509 csau_1509_i146(A[662450:660942],A[663959:662451],A[665468:663960],tree_1[442136:440628],tree_1[443645:442137]);
csa_1509 csau_1509_i147(A[666977:665469],A[668486:666978],A[669995:668487],tree_1[445154:443646],tree_1[446663:445155]);
csa_1509 csau_1509_i148(A[671504:669996],A[673013:671505],A[674522:673014],tree_1[448172:446664],tree_1[449681:448173]);
csa_1509 csau_1509_i149(A[676031:674523],A[677540:676032],A[679049:677541],tree_1[451190:449682],tree_1[452699:451191]);
csa_1509 csau_1509_i150(A[680558:679050],A[682067:680559],A[683576:682068],tree_1[454208:452700],tree_1[455717:454209]);
csa_1509 csau_1509_i151(A[685085:683577],A[686594:685086],A[688103:686595],tree_1[457226:455718],tree_1[458735:457227]);
csa_1509 csau_1509_i152(A[689612:688104],A[691121:689613],A[692630:691122],tree_1[460244:458736],tree_1[461753:460245]);
csa_1509 csau_1509_i153(A[694139:692631],A[695648:694140],A[697157:695649],tree_1[463262:461754],tree_1[464771:463263]);
csa_1509 csau_1509_i154(A[698666:697158],A[700175:698667],A[701684:700176],tree_1[466280:464772],tree_1[467789:466281]);
csa_1509 csau_1509_i155(A[703193:701685],A[704702:703194],A[706211:704703],tree_1[469298:467790],tree_1[470807:469299]);
csa_1509 csau_1509_i156(A[707720:706212],A[709229:707721],A[710738:709230],tree_1[472316:470808],tree_1[473825:472317]);
csa_1509 csau_1509_i157(A[712247:710739],A[713756:712248],A[715265:713757],tree_1[475334:473826],tree_1[476843:475335]);
csa_1509 csau_1509_i158(A[716774:715266],A[718283:716775],A[719792:718284],tree_1[478352:476844],tree_1[479861:478353]);
csa_1509 csau_1509_i159(A[721301:719793],A[722810:721302],A[724319:722811],tree_1[481370:479862],tree_1[482879:481371]);
csa_1509 csau_1509_i160(A[725828:724320],A[727337:725829],A[728846:727338],tree_1[484388:482880],tree_1[485897:484389]);
csa_1509 csau_1509_i161(A[730355:728847],A[731864:730356],A[733373:731865],tree_1[487406:485898],tree_1[488915:487407]);
csa_1509 csau_1509_i162(A[734882:733374],A[736391:734883],A[737900:736392],tree_1[490424:488916],tree_1[491933:490425]);
csa_1509 csau_1509_i163(A[739409:737901],A[740918:739410],A[742427:740919],tree_1[493442:491934],tree_1[494951:493443]);
csa_1509 csau_1509_i164(A[743936:742428],A[745445:743937],A[746954:745446],tree_1[496460:494952],tree_1[497969:496461]);
csa_1509 csau_1509_i165(A[748463:746955],A[749972:748464],A[751481:749973],tree_1[499478:497970],tree_1[500987:499479]);
csa_1509 csau_1509_i166(A[752990:751482],A[754499:752991],A[756008:754500],tree_1[502496:500988],tree_1[504005:502497]);
csa_1509 csau_1509_i167(A[757517:756009],A[759026:757518],A[760535:759027],tree_1[505514:504006],tree_1[507023:505515]);
csa_1509 csau_1509_i168(A[762044:760536],A[763553:762045],A[765062:763554],tree_1[508532:507024],tree_1[510041:508533]);
csa_1509 csau_1509_i169(A[766571:765063],A[768080:766572],A[769589:768081],tree_1[511550:510042],tree_1[513059:511551]);
csa_1509 csau_1509_i170(A[771098:769590],A[772607:771099],A[774116:772608],tree_1[514568:513060],tree_1[516077:514569]);
csa_1509 csau_1509_i171(A[775625:774117],A[777134:775626],A[778643:777135],tree_1[517586:516078],tree_1[519095:517587]);
csa_1509 csau_1509_i172(A[780152:778644],A[781661:780153],A[783170:781662],tree_1[520604:519096],tree_1[522113:520605]);
csa_1509 csau_1509_i173(A[784679:783171],A[786188:784680],A[787697:786189],tree_1[523622:522114],tree_1[525131:523623]);
csa_1509 csau_1509_i174(A[789206:787698],A[790715:789207],A[792224:790716],tree_1[526640:525132],tree_1[528149:526641]);
csa_1509 csau_1509_i175(A[793733:792225],A[795242:793734],A[796751:795243],tree_1[529658:528150],tree_1[531167:529659]);
csa_1509 csau_1509_i176(A[798260:796752],A[799769:798261],A[801278:799770],tree_1[532676:531168],tree_1[534185:532677]);
csa_1509 csau_1509_i177(A[802787:801279],A[804296:802788],A[805805:804297],tree_1[535694:534186],tree_1[537203:535695]);
csa_1509 csau_1509_i178(A[807314:805806],A[808823:807315],A[810332:808824],tree_1[538712:537204],tree_1[540221:538713]);
csa_1509 csau_1509_i179(A[811841:810333],A[813350:811842],A[814859:813351],tree_1[541730:540222],tree_1[543239:541731]);
csa_1509 csau_1509_i180(A[816368:814860],A[817877:816369],A[819386:817878],tree_1[544748:543240],tree_1[546257:544749]);
csa_1509 csau_1509_i181(A[820895:819387],A[822404:820896],A[823913:822405],tree_1[547766:546258],tree_1[549275:547767]);
csa_1509 csau_1509_i182(A[825422:823914],A[826931:825423],A[828440:826932],tree_1[550784:549276],tree_1[552293:550785]);
csa_1509 csau_1509_i183(A[829949:828441],A[831458:829950],A[832967:831459],tree_1[553802:552294],tree_1[555311:553803]);
csa_1509 csau_1509_i184(A[834476:832968],A[835985:834477],A[837494:835986],tree_1[556820:555312],tree_1[558329:556821]);
csa_1509 csau_1509_i185(A[839003:837495],A[840512:839004],A[842021:840513],tree_1[559838:558330],tree_1[561347:559839]);
csa_1509 csau_1509_i186(A[843530:842022],A[845039:843531],A[846548:845040],tree_1[562856:561348],tree_1[564365:562857]);
csa_1509 csau_1509_i187(A[848057:846549],A[849566:848058],A[851075:849567],tree_1[565874:564366],tree_1[567383:565875]);
csa_1509 csau_1509_i188(A[852584:851076],A[854093:852585],A[855602:854094],tree_1[568892:567384],tree_1[570401:568893]);
csa_1509 csau_1509_i189(A[857111:855603],A[858620:857112],A[860129:858621],tree_1[571910:570402],tree_1[573419:571911]);
csa_1509 csau_1509_i190(A[861638:860130],A[863147:861639],A[864656:863148],tree_1[574928:573420],tree_1[576437:574929]);
csa_1509 csau_1509_i191(A[866165:864657],A[867674:866166],A[869183:867675],tree_1[577946:576438],tree_1[579455:577947]);
csa_1509 csau_1509_i192(A[870692:869184],A[872201:870693],A[873710:872202],tree_1[580964:579456],tree_1[582473:580965]);
csa_1509 csau_1509_i193(A[875219:873711],A[876728:875220],A[878237:876729],tree_1[583982:582474],tree_1[585491:583983]);
csa_1509 csau_1509_i194(A[879746:878238],A[881255:879747],A[882764:881256],tree_1[587000:585492],tree_1[588509:587001]);
csa_1509 csau_1509_i195(A[884273:882765],A[885782:884274],A[887291:885783],tree_1[590018:588510],tree_1[591527:590019]);
csa_1509 csau_1509_i196(A[888800:887292],A[890309:888801],A[891818:890310],tree_1[593036:591528],tree_1[594545:593037]);
csa_1509 csau_1509_i197(A[893327:891819],A[894836:893328],A[896345:894837],tree_1[596054:594546],tree_1[597563:596055]);
csa_1509 csau_1509_i198(A[897854:896346],A[899363:897855],A[900872:899364],tree_1[599072:597564],tree_1[600581:599073]);
csa_1509 csau_1509_i199(A[902381:900873],A[903890:902382],A[905399:903891],tree_1[602090:600582],tree_1[603599:602091]);
csa_1509 csau_1509_i200(A[906908:905400],A[908417:906909],A[909926:908418],tree_1[605108:603600],tree_1[606617:605109]);
csa_1509 csau_1509_i201(A[911435:909927],A[912944:911436],A[914453:912945],tree_1[608126:606618],tree_1[609635:608127]);
csa_1509 csau_1509_i202(A[915962:914454],A[917471:915963],A[918980:917472],tree_1[611144:609636],tree_1[612653:611145]);
csa_1509 csau_1509_i203(A[920489:918981],A[921998:920490],A[923507:921999],tree_1[614162:612654],tree_1[615671:614163]);
csa_1509 csau_1509_i204(A[925016:923508],A[926525:925017],A[928034:926526],tree_1[617180:615672],tree_1[618689:617181]);
csa_1509 csau_1509_i205(A[929543:928035],A[931052:929544],A[932561:931053],tree_1[620198:618690],tree_1[621707:620199]);
csa_1509 csau_1509_i206(A[934070:932562],A[935579:934071],A[937088:935580],tree_1[623216:621708],tree_1[624725:623217]);
csa_1509 csau_1509_i207(A[938597:937089],A[940106:938598],A[941615:940107],tree_1[626234:624726],tree_1[627743:626235]);
csa_1509 csau_1509_i208(A[943124:941616],A[944633:943125],A[946142:944634],tree_1[629252:627744],tree_1[630761:629253]);
csa_1509 csau_1509_i209(A[947651:946143],A[949160:947652],A[950669:949161],tree_1[632270:630762],tree_1[633779:632271]);
csa_1509 csau_1509_i210(A[952178:950670],A[953687:952179],A[955196:953688],tree_1[635288:633780],tree_1[636797:635289]);
csa_1509 csau_1509_i211(A[956705:955197],A[958214:956706],A[959723:958215],tree_1[638306:636798],tree_1[639815:638307]);
csa_1509 csau_1509_i212(A[961232:959724],A[962741:961233],A[964250:962742],tree_1[641324:639816],tree_1[642833:641325]);
csa_1509 csau_1509_i213(A[965759:964251],A[967268:965760],A[968777:967269],tree_1[644342:642834],tree_1[645851:644343]);
csa_1509 csau_1509_i214(A[970286:968778],A[971795:970287],A[973304:971796],tree_1[647360:645852],tree_1[648869:647361]);
csa_1509 csau_1509_i215(A[974813:973305],A[976322:974814],A[977831:976323],tree_1[650378:648870],tree_1[651887:650379]);
csa_1509 csau_1509_i216(A[979340:977832],A[980849:979341],A[982358:980850],tree_1[653396:651888],tree_1[654905:653397]);
csa_1509 csau_1509_i217(A[983867:982359],A[985376:983868],A[986885:985377],tree_1[656414:654906],tree_1[657923:656415]);
csa_1509 csau_1509_i218(A[988394:986886],A[989903:988395],A[991412:989904],tree_1[659432:657924],tree_1[660941:659433]);
csa_1509 csau_1509_i219(A[992921:991413],A[994430:992922],A[995939:994431],tree_1[662450:660942],tree_1[663959:662451]);
csa_1509 csau_1509_i220(A[997448:995940],A[998957:997449],A[1000466:998958],tree_1[665468:663960],tree_1[666977:665469]);
csa_1509 csau_1509_i221(A[1001975:1000467],A[1003484:1001976],A[1004993:1003485],tree_1[668486:666978],tree_1[669995:668487]);
csa_1509 csau_1509_i222(A[1006502:1004994],A[1008011:1006503],A[1009520:1008012],tree_1[671504:669996],tree_1[673013:671505]);
csa_1509 csau_1509_i223(A[1011029:1009521],A[1012538:1011030],A[1014047:1012539],tree_1[674522:673014],tree_1[676031:674523]);
csa_1509 csau_1509_i224(A[1015556:1014048],A[1017065:1015557],A[1018574:1017066],tree_1[677540:676032],tree_1[679049:677541]);
csa_1509 csau_1509_i225(A[1020083:1018575],A[1021592:1020084],A[1023101:1021593],tree_1[680558:679050],tree_1[682067:680559]);
csa_1509 csau_1509_i226(A[1024610:1023102],A[1026119:1024611],A[1027628:1026120],tree_1[683576:682068],tree_1[685085:683577]);
csa_1509 csau_1509_i227(A[1029137:1027629],A[1030646:1029138],A[1032155:1030647],tree_1[686594:685086],tree_1[688103:686595]);
csa_1509 csau_1509_i228(A[1033664:1032156],A[1035173:1033665],A[1036682:1035174],tree_1[689612:688104],tree_1[691121:689613]);
csa_1509 csau_1509_i229(A[1038191:1036683],A[1039700:1038192],A[1041209:1039701],tree_1[692630:691122],tree_1[694139:692631]);
csa_1509 csau_1509_i230(A[1042718:1041210],A[1044227:1042719],A[1045736:1044228],tree_1[695648:694140],tree_1[697157:695649]);
csa_1509 csau_1509_i231(A[1047245:1045737],A[1048754:1047246],A[1050263:1048755],tree_1[698666:697158],tree_1[700175:698667]);
csa_1509 csau_1509_i232(A[1051772:1050264],A[1053281:1051773],A[1054790:1053282],tree_1[701684:700176],tree_1[703193:701685]);
csa_1509 csau_1509_i233(A[1056299:1054791],A[1057808:1056300],A[1059317:1057809],tree_1[704702:703194],tree_1[706211:704703]);
csa_1509 csau_1509_i234(A[1060826:1059318],A[1062335:1060827],A[1063844:1062336],tree_1[707720:706212],tree_1[709229:707721]);
csa_1509 csau_1509_i235(A[1065353:1063845],A[1066862:1065354],A[1068371:1066863],tree_1[710738:709230],tree_1[712247:710739]);
csa_1509 csau_1509_i236(A[1069880:1068372],A[1071389:1069881],A[1072898:1071390],tree_1[713756:712248],tree_1[715265:713757]);
csa_1509 csau_1509_i237(A[1074407:1072899],A[1075916:1074408],A[1077425:1075917],tree_1[716774:715266],tree_1[718283:716775]);
csa_1509 csau_1509_i238(A[1078934:1077426],A[1080443:1078935],A[1081952:1080444],tree_1[719792:718284],tree_1[721301:719793]);
csa_1509 csau_1509_i239(A[1083461:1081953],A[1084970:1083462],A[1086479:1084971],tree_1[722810:721302],tree_1[724319:722811]);
csa_1509 csau_1509_i240(A[1087988:1086480],A[1089497:1087989],A[1091006:1089498],tree_1[725828:724320],tree_1[727337:725829]);
csa_1509 csau_1509_i241(A[1092515:1091007],A[1094024:1092516],A[1095533:1094025],tree_1[728846:727338],tree_1[730355:728847]);
csa_1509 csau_1509_i242(A[1097042:1095534],A[1098551:1097043],A[1100060:1098552],tree_1[731864:730356],tree_1[733373:731865]);
csa_1509 csau_1509_i243(A[1101569:1100061],A[1103078:1101570],A[1104587:1103079],tree_1[734882:733374],tree_1[736391:734883]);
csa_1509 csau_1509_i244(A[1106096:1104588],A[1107605:1106097],A[1109114:1107606],tree_1[737900:736392],tree_1[739409:737901]);
csa_1509 csau_1509_i245(A[1110623:1109115],A[1112132:1110624],A[1113641:1112133],tree_1[740918:739410],tree_1[742427:740919]);
csa_1509 csau_1509_i246(A[1115150:1113642],A[1116659:1115151],A[1118168:1116660],tree_1[743936:742428],tree_1[745445:743937]);
csa_1509 csau_1509_i247(A[1119677:1118169],A[1121186:1119678],A[1122695:1121187],tree_1[746954:745446],tree_1[748463:746955]);
csa_1509 csau_1509_i248(A[1124204:1122696],A[1125713:1124205],A[1127222:1125714],tree_1[749972:748464],tree_1[751481:749973]);
csa_1509 csau_1509_i249(A[1128731:1127223],A[1130240:1128732],A[1131749:1130241],tree_1[752990:751482],tree_1[754499:752991]);
csa_1509 csau_1509_i250(A[1133258:1131750],A[1134767:1133259],A[1136276:1134768],tree_1[756008:754500],tree_1[757517:756009]);
csa_1509 csau_1509_i251(A[1137785:1136277],A[1139294:1137786],A[1140803:1139295],tree_1[759026:757518],tree_1[760535:759027]);
csa_1509 csau_1509_i252(A[1142312:1140804],A[1143821:1142313],A[1145330:1143822],tree_1[762044:760536],tree_1[763553:762045]);
csa_1509 csau_1509_i253(A[1146839:1145331],A[1148348:1146840],A[1149857:1148349],tree_1[765062:763554],tree_1[766571:765063]);
csa_1509 csau_1509_i254(A[1151366:1149858],A[1152875:1151367],A[1154384:1152876],tree_1[768080:766572],tree_1[769589:768081]);
csa_1509 csau_1509_i255(A[1155893:1154385],A[1157402:1155894],A[1158911:1157403],tree_1[771098:769590],tree_1[772607:771099]);
csa_1509 csau_1509_i256(A[1160420:1158912],A[1161929:1160421],A[1163438:1161930],tree_1[774116:772608],tree_1[775625:774117]);
csa_1509 csau_1509_i257(A[1164947:1163439],A[1166456:1164948],A[1167965:1166457],tree_1[777134:775626],tree_1[778643:777135]);
csa_1509 csau_1509_i258(A[1169474:1167966],A[1170983:1169475],A[1172492:1170984],tree_1[780152:778644],tree_1[781661:780153]);
csa_1509 csau_1509_i259(A[1174001:1172493],A[1175510:1174002],A[1177019:1175511],tree_1[783170:781662],tree_1[784679:783171]);
csa_1509 csau_1509_i260(A[1178528:1177020],A[1180037:1178529],A[1181546:1180038],tree_1[786188:784680],tree_1[787697:786189]);
csa_1509 csau_1509_i261(A[1183055:1181547],A[1184564:1183056],A[1186073:1184565],tree_1[789206:787698],tree_1[790715:789207]);
csa_1509 csau_1509_i262(A[1187582:1186074],A[1189091:1187583],A[1190600:1189092],tree_1[792224:790716],tree_1[793733:792225]);
csa_1509 csau_1509_i263(A[1192109:1190601],A[1193618:1192110],A[1195127:1193619],tree_1[795242:793734],tree_1[796751:795243]);
csa_1509 csau_1509_i264(A[1196636:1195128],A[1198145:1196637],A[1199654:1198146],tree_1[798260:796752],tree_1[799769:798261]);
csa_1509 csau_1509_i265(A[1201163:1199655],A[1202672:1201164],A[1204181:1202673],tree_1[801278:799770],tree_1[802787:801279]);
csa_1509 csau_1509_i266(A[1205690:1204182],A[1207199:1205691],A[1208708:1207200],tree_1[804296:802788],tree_1[805805:804297]);
csa_1509 csau_1509_i267(A[1210217:1208709],A[1211726:1210218],A[1213235:1211727],tree_1[807314:805806],tree_1[808823:807315]);
csa_1509 csau_1509_i268(A[1214744:1213236],A[1216253:1214745],A[1217762:1216254],tree_1[810332:808824],tree_1[811841:810333]);
csa_1509 csau_1509_i269(A[1219271:1217763],A[1220780:1219272],A[1222289:1220781],tree_1[813350:811842],tree_1[814859:813351]);
csa_1509 csau_1509_i270(A[1223798:1222290],A[1225307:1223799],A[1226816:1225308],tree_1[816368:814860],tree_1[817877:816369]);
csa_1509 csau_1509_i271(A[1228325:1226817],A[1229834:1228326],A[1231343:1229835],tree_1[819386:817878],tree_1[820895:819387]);
csa_1509 csau_1509_i272(A[1232852:1231344],A[1234361:1232853],A[1235870:1234362],tree_1[822404:820896],tree_1[823913:822405]);
csa_1509 csau_1509_i273(A[1237379:1235871],A[1238888:1237380],A[1240397:1238889],tree_1[825422:823914],tree_1[826931:825423]);
csa_1509 csau_1509_i274(A[1241906:1240398],A[1243415:1241907],A[1244924:1243416],tree_1[828440:826932],tree_1[829949:828441]);
csa_1509 csau_1509_i275(A[1246433:1244925],A[1247942:1246434],A[1249451:1247943],tree_1[831458:829950],tree_1[832967:831459]);
csa_1509 csau_1509_i276(A[1250960:1249452],A[1252469:1250961],A[1253978:1252470],tree_1[834476:832968],tree_1[835985:834477]);
csa_1509 csau_1509_i277(A[1255487:1253979],A[1256996:1255488],A[1258505:1256997],tree_1[837494:835986],tree_1[839003:837495]);
csa_1509 csau_1509_i278(A[1260014:1258506],A[1261523:1260015],A[1263032:1261524],tree_1[840512:839004],tree_1[842021:840513]);
csa_1509 csau_1509_i279(A[1264541:1263033],A[1266050:1264542],A[1267559:1266051],tree_1[843530:842022],tree_1[845039:843531]);
csa_1509 csau_1509_i280(A[1269068:1267560],A[1270577:1269069],A[1272086:1270578],tree_1[846548:845040],tree_1[848057:846549]);
csa_1509 csau_1509_i281(A[1273595:1272087],A[1275104:1273596],A[1276613:1275105],tree_1[849566:848058],tree_1[851075:849567]);
csa_1509 csau_1509_i282(A[1278122:1276614],A[1279631:1278123],A[1281140:1279632],tree_1[852584:851076],tree_1[854093:852585]);
csa_1509 csau_1509_i283(A[1282649:1281141],A[1284158:1282650],A[1285667:1284159],tree_1[855602:854094],tree_1[857111:855603]);
csa_1509 csau_1509_i284(A[1287176:1285668],A[1288685:1287177],A[1290194:1288686],tree_1[858620:857112],tree_1[860129:858621]);
csa_1509 csau_1509_i285(A[1291703:1290195],A[1293212:1291704],A[1294721:1293213],tree_1[861638:860130],tree_1[863147:861639]);
csa_1509 csau_1509_i286(A[1296230:1294722],A[1297739:1296231],A[1299248:1297740],tree_1[864656:863148],tree_1[866165:864657]);
csa_1509 csau_1509_i287(A[1300757:1299249],A[1302266:1300758],A[1303775:1302267],tree_1[867674:866166],tree_1[869183:867675]);
csa_1509 csau_1509_i288(A[1305284:1303776],A[1306793:1305285],A[1308302:1306794],tree_1[870692:869184],tree_1[872201:870693]);
csa_1509 csau_1509_i289(A[1309811:1308303],A[1311320:1309812],A[1312829:1311321],tree_1[873710:872202],tree_1[875219:873711]);
csa_1509 csau_1509_i290(A[1314338:1312830],A[1315847:1314339],A[1317356:1315848],tree_1[876728:875220],tree_1[878237:876729]);
csa_1509 csau_1509_i291(A[1318865:1317357],A[1320374:1318866],A[1321883:1320375],tree_1[879746:878238],tree_1[881255:879747]);
csa_1509 csau_1509_i292(A[1323392:1321884],A[1324901:1323393],A[1326410:1324902],tree_1[882764:881256],tree_1[884273:882765]);
csa_1509 csau_1509_i293(A[1327919:1326411],A[1329428:1327920],A[1330937:1329429],tree_1[885782:884274],tree_1[887291:885783]);
csa_1509 csau_1509_i294(A[1332446:1330938],A[1333955:1332447],A[1335464:1333956],tree_1[888800:887292],tree_1[890309:888801]);
csa_1509 csau_1509_i295(A[1336973:1335465],A[1338482:1336974],A[1339991:1338483],tree_1[891818:890310],tree_1[893327:891819]);
csa_1509 csau_1509_i296(A[1341500:1339992],A[1343009:1341501],A[1344518:1343010],tree_1[894836:893328],tree_1[896345:894837]);
csa_1509 csau_1509_i297(A[1346027:1344519],A[1347536:1346028],A[1349045:1347537],tree_1[897854:896346],tree_1[899363:897855]);
csa_1509 csau_1509_i298(A[1350554:1349046],A[1352063:1350555],A[1353572:1352064],tree_1[900872:899364],tree_1[902381:900873]);
csa_1509 csau_1509_i299(A[1355081:1353573],A[1356590:1355082],A[1358099:1356591],tree_1[903890:902382],tree_1[905399:903891]);
csa_1509 csau_1509_i300(A[1359608:1358100],A[1361117:1359609],A[1362626:1361118],tree_1[906908:905400],tree_1[908417:906909]);
csa_1509 csau_1509_i301(A[1364135:1362627],A[1365644:1364136],A[1367153:1365645],tree_1[909926:908418],tree_1[911435:909927]);
csa_1509 csau_1509_i302(A[1368662:1367154],A[1370171:1368663],A[1371680:1370172],tree_1[912944:911436],tree_1[914453:912945]);
csa_1509 csau_1509_i303(A[1373189:1371681],A[1374698:1373190],A[1376207:1374699],tree_1[915962:914454],tree_1[917471:915963]);
csa_1509 csau_1509_i304(A[1377716:1376208],A[1379225:1377717],A[1380734:1379226],tree_1[918980:917472],tree_1[920489:918981]);
csa_1509 csau_1509_i305(A[1382243:1380735],A[1383752:1382244],A[1385261:1383753],tree_1[921998:920490],tree_1[923507:921999]);
csa_1509 csau_1509_i306(A[1386770:1385262],A[1388279:1386771],A[1389788:1388280],tree_1[925016:923508],tree_1[926525:925017]);
csa_1509 csau_1509_i307(A[1391297:1389789],A[1392806:1391298],A[1394315:1392807],tree_1[928034:926526],tree_1[929543:928035]);
csa_1509 csau_1509_i308(A[1395824:1394316],A[1397333:1395825],A[1398842:1397334],tree_1[931052:929544],tree_1[932561:931053]);
csa_1509 csau_1509_i309(A[1400351:1398843],A[1401860:1400352],A[1403369:1401861],tree_1[934070:932562],tree_1[935579:934071]);
csa_1509 csau_1509_i310(A[1404878:1403370],A[1406387:1404879],A[1407896:1406388],tree_1[937088:935580],tree_1[938597:937089]);
csa_1509 csau_1509_i311(A[1409405:1407897],A[1410914:1409406],A[1412423:1410915],tree_1[940106:938598],tree_1[941615:940107]);
csa_1509 csau_1509_i312(A[1413932:1412424],A[1415441:1413933],A[1416950:1415442],tree_1[943124:941616],tree_1[944633:943125]);
csa_1509 csau_1509_i313(A[1418459:1416951],A[1419968:1418460],A[1421477:1419969],tree_1[946142:944634],tree_1[947651:946143]);
csa_1509 csau_1509_i314(A[1422986:1421478],A[1424495:1422987],A[1426004:1424496],tree_1[949160:947652],tree_1[950669:949161]);
csa_1509 csau_1509_i315(A[1427513:1426005],A[1429022:1427514],A[1430531:1429023],tree_1[952178:950670],tree_1[953687:952179]);
csa_1509 csau_1509_i316(A[1432040:1430532],A[1433549:1432041],A[1435058:1433550],tree_1[955196:953688],tree_1[956705:955197]);
csa_1509 csau_1509_i317(A[1436567:1435059],A[1438076:1436568],A[1439585:1438077],tree_1[958214:956706],tree_1[959723:958215]);
csa_1509 csau_1509_i318(A[1441094:1439586],A[1442603:1441095],A[1444112:1442604],tree_1[961232:959724],tree_1[962741:961233]);
csa_1509 csau_1509_i319(A[1445621:1444113],A[1447130:1445622],A[1448639:1447131],tree_1[964250:962742],tree_1[965759:964251]);
csa_1509 csau_1509_i320(A[1450148:1448640],A[1451657:1450149],A[1453166:1451658],tree_1[967268:965760],tree_1[968777:967269]);
csa_1509 csau_1509_i321(A[1454675:1453167],A[1456184:1454676],A[1457693:1456185],tree_1[970286:968778],tree_1[971795:970287]);
csa_1509 csau_1509_i322(A[1459202:1457694],A[1460711:1459203],A[1462220:1460712],tree_1[973304:971796],tree_1[974813:973305]);
csa_1509 csau_1509_i323(A[1463729:1462221],A[1465238:1463730],A[1466747:1465239],tree_1[976322:974814],tree_1[977831:976323]);
csa_1509 csau_1509_i324(A[1468256:1466748],A[1469765:1468257],A[1471274:1469766],tree_1[979340:977832],tree_1[980849:979341]);
csa_1509 csau_1509_i325(A[1472783:1471275],A[1474292:1472784],A[1475801:1474293],tree_1[982358:980850],tree_1[983867:982359]);
csa_1509 csau_1509_i326(A[1477310:1475802],A[1478819:1477311],A[1480328:1478820],tree_1[985376:983868],tree_1[986885:985377]);
csa_1509 csau_1509_i327(A[1481837:1480329],A[1483346:1481838],A[1484855:1483347],tree_1[988394:986886],tree_1[989903:988395]);
csa_1509 csau_1509_i328(A[1486364:1484856],A[1487873:1486365],A[1489382:1487874],tree_1[991412:989904],tree_1[992921:991413]);
csa_1509 csau_1509_i329(A[1490891:1489383],A[1492400:1490892],A[1493909:1492401],tree_1[994430:992922],tree_1[995939:994431]);
csa_1509 csau_1509_i330(A[1495418:1493910],A[1496927:1495419],A[1498436:1496928],tree_1[997448:995940],tree_1[998957:997449]);
csa_1509 csau_1509_i331(A[1499945:1498437],A[1501454:1499946],A[1502963:1501455],tree_1[1000466:998958],tree_1[1001975:1000467]);
csa_1509 csau_1509_i332(A[1504472:1502964],A[1505981:1504473],A[1507490:1505982],tree_1[1003484:1001976],tree_1[1004993:1003485]);
csa_1509 csau_1509_i333(A[1508999:1507491],A[1510508:1509000],A[1512017:1510509],tree_1[1006502:1004994],tree_1[1008011:1006503]);
csa_1509 csau_1509_i334(A[1513526:1512018],A[1515035:1513527],A[1516544:1515036],tree_1[1009520:1008012],tree_1[1011029:1009521]);
csa_1509 csau_1509_i335(A[1518053:1516545],A[1519562:1518054],A[1521071:1519563],tree_1[1012538:1011030],tree_1[1014047:1012539]);
csa_1509 csau_1509_i336(A[1522580:1521072],A[1524089:1522581],A[1525598:1524090],tree_1[1015556:1014048],tree_1[1017065:1015557]);
csa_1509 csau_1509_i337(A[1527107:1525599],A[1528616:1527108],A[1530125:1528617],tree_1[1018574:1017066],tree_1[1020083:1018575]);
csa_1509 csau_1509_i338(A[1531634:1530126],A[1533143:1531635],A[1534652:1533144],tree_1[1021592:1020084],tree_1[1023101:1021593]);
csa_1509 csau_1509_i339(A[1536161:1534653],A[1537670:1536162],A[1539179:1537671],tree_1[1024610:1023102],tree_1[1026119:1024611]);
csa_1509 csau_1509_i340(A[1540688:1539180],A[1542197:1540689],A[1543706:1542198],tree_1[1027628:1026120],tree_1[1029137:1027629]);
csa_1509 csau_1509_i341(A[1545215:1543707],A[1546724:1545216],A[1548233:1546725],tree_1[1030646:1029138],tree_1[1032155:1030647]);
csa_1509 csau_1509_i342(A[1549742:1548234],A[1551251:1549743],A[1552760:1551252],tree_1[1033664:1032156],tree_1[1035173:1033665]);
csa_1509 csau_1509_i343(A[1554269:1552761],A[1555778:1554270],A[1557287:1555779],tree_1[1036682:1035174],tree_1[1038191:1036683]);
csa_1509 csau_1509_i344(A[1558796:1557288],A[1560305:1558797],A[1561814:1560306],tree_1[1039700:1038192],tree_1[1041209:1039701]);
csa_1509 csau_1509_i345(A[1563323:1561815],A[1564832:1563324],A[1566341:1564833],tree_1[1042718:1041210],tree_1[1044227:1042719]);
csa_1509 csau_1509_i346(A[1567850:1566342],A[1569359:1567851],A[1570868:1569360],tree_1[1045736:1044228],tree_1[1047245:1045737]);
csa_1509 csau_1509_i347(A[1572377:1570869],A[1573886:1572378],A[1575395:1573887],tree_1[1048754:1047246],tree_1[1050263:1048755]);
csa_1509 csau_1509_i348(A[1576904:1575396],A[1578413:1576905],A[1579922:1578414],tree_1[1051772:1050264],tree_1[1053281:1051773]);
csa_1509 csau_1509_i349(A[1581431:1579923],A[1582940:1581432],A[1584449:1582941],tree_1[1054790:1053282],tree_1[1056299:1054791]);
csa_1509 csau_1509_i350(A[1585958:1584450],A[1587467:1585959],A[1588976:1587468],tree_1[1057808:1056300],tree_1[1059317:1057809]);
csa_1509 csau_1509_i351(A[1590485:1588977],A[1591994:1590486],A[1593503:1591995],tree_1[1060826:1059318],tree_1[1062335:1060827]);
csa_1509 csau_1509_i352(A[1595012:1593504],A[1596521:1595013],A[1598030:1596522],tree_1[1063844:1062336],tree_1[1065353:1063845]);
csa_1509 csau_1509_i353(A[1599539:1598031],A[1601048:1599540],A[1602557:1601049],tree_1[1066862:1065354],tree_1[1068371:1066863]);
csa_1509 csau_1509_i354(A[1604066:1602558],A[1605575:1604067],A[1607084:1605576],tree_1[1069880:1068372],tree_1[1071389:1069881]);
csa_1509 csau_1509_i355(A[1608593:1607085],A[1610102:1608594],A[1611611:1610103],tree_1[1072898:1071390],tree_1[1074407:1072899]);
csa_1509 csau_1509_i356(A[1613120:1611612],A[1614629:1613121],A[1616138:1614630],tree_1[1075916:1074408],tree_1[1077425:1075917]);
csa_1509 csau_1509_i357(A[1617647:1616139],A[1619156:1617648],A[1620665:1619157],tree_1[1078934:1077426],tree_1[1080443:1078935]);
csa_1509 csau_1509_i358(A[1622174:1620666],A[1623683:1622175],A[1625192:1623684],tree_1[1081952:1080444],tree_1[1083461:1081953]);
csa_1509 csau_1509_i359(A[1626701:1625193],A[1628210:1626702],A[1629719:1628211],tree_1[1084970:1083462],tree_1[1086479:1084971]);
csa_1509 csau_1509_i360(A[1631228:1629720],A[1632737:1631229],A[1634246:1632738],tree_1[1087988:1086480],tree_1[1089497:1087989]);
csa_1509 csau_1509_i361(A[1635755:1634247],A[1637264:1635756],A[1638773:1637265],tree_1[1091006:1089498],tree_1[1092515:1091007]);
csa_1509 csau_1509_i362(A[1640282:1638774],A[1641791:1640283],A[1643300:1641792],tree_1[1094024:1092516],tree_1[1095533:1094025]);
csa_1509 csau_1509_i363(A[1644809:1643301],A[1646318:1644810],A[1647827:1646319],tree_1[1097042:1095534],tree_1[1098551:1097043]);
csa_1509 csau_1509_i364(A[1649336:1647828],A[1650845:1649337],A[1652354:1650846],tree_1[1100060:1098552],tree_1[1101569:1100061]);
csa_1509 csau_1509_i365(A[1653863:1652355],A[1655372:1653864],A[1656881:1655373],tree_1[1103078:1101570],tree_1[1104587:1103079]);
csa_1509 csau_1509_i366(A[1658390:1656882],A[1659899:1658391],A[1661408:1659900],tree_1[1106096:1104588],tree_1[1107605:1106097]);
csa_1509 csau_1509_i367(A[1662917:1661409],A[1664426:1662918],A[1665935:1664427],tree_1[1109114:1107606],tree_1[1110623:1109115]);
csa_1509 csau_1509_i368(A[1667444:1665936],A[1668953:1667445],A[1670462:1668954],tree_1[1112132:1110624],tree_1[1113641:1112133]);
csa_1509 csau_1509_i369(A[1671971:1670463],A[1673480:1671972],A[1674989:1673481],tree_1[1115150:1113642],tree_1[1116659:1115151]);
csa_1509 csau_1509_i370(A[1676498:1674990],A[1678007:1676499],A[1679516:1678008],tree_1[1118168:1116660],tree_1[1119677:1118169]);
csa_1509 csau_1509_i371(A[1681025:1679517],A[1682534:1681026],A[1684043:1682535],tree_1[1121186:1119678],tree_1[1122695:1121187]);
csa_1509 csau_1509_i372(A[1685552:1684044],A[1687061:1685553],A[1688570:1687062],tree_1[1124204:1122696],tree_1[1125713:1124205]);
csa_1509 csau_1509_i373(A[1690079:1688571],A[1691588:1690080],A[1693097:1691589],tree_1[1127222:1125714],tree_1[1128731:1127223]);
csa_1509 csau_1509_i374(A[1694606:1693098],A[1696115:1694607],A[1697624:1696116],tree_1[1130240:1128732],tree_1[1131749:1130241]);
csa_1509 csau_1509_i375(A[1699133:1697625],A[1700642:1699134],A[1702151:1700643],tree_1[1133258:1131750],tree_1[1134767:1133259]);
csa_1509 csau_1509_i376(A[1703660:1702152],A[1705169:1703661],A[1706678:1705170],tree_1[1136276:1134768],tree_1[1137785:1136277]);
csa_1509 csau_1509_i377(A[1708187:1706679],A[1709696:1708188],A[1711205:1709697],tree_1[1139294:1137786],tree_1[1140803:1139295]);
csa_1509 csau_1509_i378(A[1712714:1711206],A[1714223:1712715],A[1715732:1714224],tree_1[1142312:1140804],tree_1[1143821:1142313]);
csa_1509 csau_1509_i379(A[1717241:1715733],A[1718750:1717242],A[1720259:1718751],tree_1[1145330:1143822],tree_1[1146839:1145331]);
csa_1509 csau_1509_i380(A[1721768:1720260],A[1723277:1721769],A[1724786:1723278],tree_1[1148348:1146840],tree_1[1149857:1148349]);
csa_1509 csau_1509_i381(A[1726295:1724787],A[1727804:1726296],A[1729313:1727805],tree_1[1151366:1149858],tree_1[1152875:1151367]);
csa_1509 csau_1509_i382(A[1730822:1729314],A[1732331:1730823],A[1733840:1732332],tree_1[1154384:1152876],tree_1[1155893:1154385]);
csa_1509 csau_1509_i383(A[1735349:1733841],A[1736858:1735350],A[1738367:1736859],tree_1[1157402:1155894],tree_1[1158911:1157403]);
csa_1509 csau_1509_i384(A[1739876:1738368],A[1741385:1739877],A[1742894:1741386],tree_1[1160420:1158912],tree_1[1161929:1160421]);
csa_1509 csau_1509_i385(A[1744403:1742895],A[1745912:1744404],A[1747421:1745913],tree_1[1163438:1161930],tree_1[1164947:1163439]);
csa_1509 csau_1509_i386(A[1748930:1747422],A[1750439:1748931],A[1751948:1750440],tree_1[1166456:1164948],tree_1[1167965:1166457]);
csa_1509 csau_1509_i387(A[1753457:1751949],A[1754966:1753458],A[1756475:1754967],tree_1[1169474:1167966],tree_1[1170983:1169475]);
csa_1509 csau_1509_i388(A[1757984:1756476],A[1759493:1757985],A[1761002:1759494],tree_1[1172492:1170984],tree_1[1174001:1172493]);
csa_1509 csau_1509_i389(A[1762511:1761003],A[1764020:1762512],A[1765529:1764021],tree_1[1175510:1174002],tree_1[1177019:1175511]);
csa_1509 csau_1509_i390(A[1767038:1765530],A[1768547:1767039],A[1770056:1768548],tree_1[1178528:1177020],tree_1[1180037:1178529]);
csa_1509 csau_1509_i391(A[1771565:1770057],A[1773074:1771566],A[1774583:1773075],tree_1[1181546:1180038],tree_1[1183055:1181547]);
csa_1509 csau_1509_i392(A[1776092:1774584],A[1777601:1776093],A[1779110:1777602],tree_1[1184564:1183056],tree_1[1186073:1184565]);
csa_1509 csau_1509_i393(A[1780619:1779111],A[1782128:1780620],A[1783637:1782129],tree_1[1187582:1186074],tree_1[1189091:1187583]);
csa_1509 csau_1509_i394(A[1785146:1783638],A[1786655:1785147],A[1788164:1786656],tree_1[1190600:1189092],tree_1[1192109:1190601]);
csa_1509 csau_1509_i395(A[1789673:1788165],A[1791182:1789674],A[1792691:1791183],tree_1[1193618:1192110],tree_1[1195127:1193619]);
csa_1509 csau_1509_i396(A[1794200:1792692],A[1795709:1794201],A[1797218:1795710],tree_1[1196636:1195128],tree_1[1198145:1196637]);
csa_1509 csau_1509_i397(A[1798727:1797219],A[1800236:1798728],A[1801745:1800237],tree_1[1199654:1198146],tree_1[1201163:1199655]);
csa_1509 csau_1509_i398(A[1803254:1801746],A[1804763:1803255],A[1806272:1804764],tree_1[1202672:1201164],tree_1[1204181:1202673]);
csa_1509 csau_1509_i399(A[1807781:1806273],A[1809290:1807782],A[1810799:1809291],tree_1[1205690:1204182],tree_1[1207199:1205691]);
csa_1509 csau_1509_i400(A[1812308:1810800],A[1813817:1812309],A[1815326:1813818],tree_1[1208708:1207200],tree_1[1210217:1208709]);
csa_1509 csau_1509_i401(A[1816835:1815327],A[1818344:1816836],A[1819853:1818345],tree_1[1211726:1210218],tree_1[1213235:1211727]);
csa_1509 csau_1509_i402(A[1821362:1819854],A[1822871:1821363],A[1824380:1822872],tree_1[1214744:1213236],tree_1[1216253:1214745]);
csa_1509 csau_1509_i403(A[1825889:1824381],A[1827398:1825890],A[1828907:1827399],tree_1[1217762:1216254],tree_1[1219271:1217763]);
csa_1509 csau_1509_i404(A[1830416:1828908],A[1831925:1830417],A[1833434:1831926],tree_1[1220780:1219272],tree_1[1222289:1220781]);
csa_1509 csau_1509_i405(A[1834943:1833435],A[1836452:1834944],A[1837961:1836453],tree_1[1223798:1222290],tree_1[1225307:1223799]);
csa_1509 csau_1509_i406(A[1839470:1837962],A[1840979:1839471],A[1842488:1840980],tree_1[1226816:1225308],tree_1[1228325:1226817]);
csa_1509 csau_1509_i407(A[1843997:1842489],A[1845506:1843998],A[1847015:1845507],tree_1[1229834:1228326],tree_1[1231343:1229835]);
csa_1509 csau_1509_i408(A[1848524:1847016],A[1850033:1848525],A[1851542:1850034],tree_1[1232852:1231344],tree_1[1234361:1232853]);
csa_1509 csau_1509_i409(A[1853051:1851543],A[1854560:1853052],A[1856069:1854561],tree_1[1235870:1234362],tree_1[1237379:1235871]);
csa_1509 csau_1509_i410(A[1857578:1856070],A[1859087:1857579],A[1860596:1859088],tree_1[1238888:1237380],tree_1[1240397:1238889]);
csa_1509 csau_1509_i411(A[1862105:1860597],A[1863614:1862106],A[1865123:1863615],tree_1[1241906:1240398],tree_1[1243415:1241907]);
csa_1509 csau_1509_i412(A[1866632:1865124],A[1868141:1866633],A[1869650:1868142],tree_1[1244924:1243416],tree_1[1246433:1244925]);
csa_1509 csau_1509_i413(A[1871159:1869651],A[1872668:1871160],A[1874177:1872669],tree_1[1247942:1246434],tree_1[1249451:1247943]);
csa_1509 csau_1509_i414(A[1875686:1874178],A[1877195:1875687],A[1878704:1877196],tree_1[1250960:1249452],tree_1[1252469:1250961]);
csa_1509 csau_1509_i415(A[1880213:1878705],A[1881722:1880214],A[1883231:1881723],tree_1[1253978:1252470],tree_1[1255487:1253979]);
csa_1509 csau_1509_i416(A[1884740:1883232],A[1886249:1884741],A[1887758:1886250],tree_1[1256996:1255488],tree_1[1258505:1256997]);
csa_1509 csau_1509_i417(A[1889267:1887759],A[1890776:1889268],A[1892285:1890777],tree_1[1260014:1258506],tree_1[1261523:1260015]);
csa_1509 csau_1509_i418(A[1893794:1892286],A[1895303:1893795],A[1896812:1895304],tree_1[1263032:1261524],tree_1[1264541:1263033]);
csa_1509 csau_1509_i419(A[1898321:1896813],A[1899830:1898322],A[1901339:1899831],tree_1[1266050:1264542],tree_1[1267559:1266051]);
csa_1509 csau_1509_i420(A[1902848:1901340],A[1904357:1902849],A[1905866:1904358],tree_1[1269068:1267560],tree_1[1270577:1269069]);
csa_1509 csau_1509_i421(A[1907375:1905867],A[1908884:1907376],A[1910393:1908885],tree_1[1272086:1270578],tree_1[1273595:1272087]);
csa_1509 csau_1509_i422(A[1911902:1910394],A[1913411:1911903],A[1914920:1913412],tree_1[1275104:1273596],tree_1[1276613:1275105]);
csa_1509 csau_1509_i423(A[1916429:1914921],A[1917938:1916430],A[1919447:1917939],tree_1[1278122:1276614],tree_1[1279631:1278123]);
csa_1509 csau_1509_i424(A[1920956:1919448],A[1922465:1920957],A[1923974:1922466],tree_1[1281140:1279632],tree_1[1282649:1281141]);
csa_1509 csau_1509_i425(A[1925483:1923975],A[1926992:1925484],A[1928501:1926993],tree_1[1284158:1282650],tree_1[1285667:1284159]);
csa_1509 csau_1509_i426(A[1930010:1928502],A[1931519:1930011],A[1933028:1931520],tree_1[1287176:1285668],tree_1[1288685:1287177]);
csa_1509 csau_1509_i427(A[1934537:1933029],A[1936046:1934538],A[1937555:1936047],tree_1[1290194:1288686],tree_1[1291703:1290195]);
csa_1509 csau_1509_i428(A[1939064:1937556],A[1940573:1939065],A[1942082:1940574],tree_1[1293212:1291704],tree_1[1294721:1293213]);
csa_1509 csau_1509_i429(A[1943591:1942083],A[1945100:1943592],A[1946609:1945101],tree_1[1296230:1294722],tree_1[1297739:1296231]);
csa_1509 csau_1509_i430(A[1948118:1946610],A[1949627:1948119],A[1951136:1949628],tree_1[1299248:1297740],tree_1[1300757:1299249]);
csa_1509 csau_1509_i431(A[1952645:1951137],A[1954154:1952646],A[1955663:1954155],tree_1[1302266:1300758],tree_1[1303775:1302267]);
csa_1509 csau_1509_i432(A[1957172:1955664],A[1958681:1957173],A[1960190:1958682],tree_1[1305284:1303776],tree_1[1306793:1305285]);
csa_1509 csau_1509_i433(A[1961699:1960191],A[1963208:1961700],A[1964717:1963209],tree_1[1308302:1306794],tree_1[1309811:1308303]);
csa_1509 csau_1509_i434(A[1966226:1964718],A[1967735:1966227],A[1969244:1967736],tree_1[1311320:1309812],tree_1[1312829:1311321]);
csa_1509 csau_1509_i435(A[1970753:1969245],A[1972262:1970754],A[1973771:1972263],tree_1[1314338:1312830],tree_1[1315847:1314339]);
csa_1509 csau_1509_i436(A[1975280:1973772],A[1976789:1975281],A[1978298:1976790],tree_1[1317356:1315848],tree_1[1318865:1317357]);
csa_1509 csau_1509_i437(A[1979807:1978299],A[1981316:1979808],A[1982825:1981317],tree_1[1320374:1318866],tree_1[1321883:1320375]);
csa_1509 csau_1509_i438(A[1984334:1982826],A[1985843:1984335],A[1987352:1985844],tree_1[1323392:1321884],tree_1[1324901:1323393]);
csa_1509 csau_1509_i439(A[1988861:1987353],A[1990370:1988862],A[1991879:1990371],tree_1[1326410:1324902],tree_1[1327919:1326411]);
csa_1509 csau_1509_i440(A[1993388:1991880],A[1994897:1993389],A[1996406:1994898],tree_1[1329428:1327920],tree_1[1330937:1329429]);
csa_1509 csau_1509_i441(A[1997915:1996407],A[1999424:1997916],A[2000933:1999425],tree_1[1332446:1330938],tree_1[1333955:1332447]);
csa_1509 csau_1509_i442(A[2002442:2000934],A[2003951:2002443],A[2005460:2003952],tree_1[1335464:1333956],tree_1[1336973:1335465]);
csa_1509 csau_1509_i443(A[2006969:2005461],A[2008478:2006970],A[2009987:2008479],tree_1[1338482:1336974],tree_1[1339991:1338483]);
csa_1509 csau_1509_i444(A[2011496:2009988],A[2013005:2011497],A[2014514:2013006],tree_1[1341500:1339992],tree_1[1343009:1341501]);
csa_1509 csau_1509_i445(A[2016023:2014515],A[2017532:2016024],A[2019041:2017533],tree_1[1344518:1343010],tree_1[1346027:1344519]);
csa_1509 csau_1509_i446(A[2020550:2019042],A[2022059:2020551],A[2023568:2022060],tree_1[1347536:1346028],tree_1[1349045:1347537]);
csa_1509 csau_1509_i447(A[2025077:2023569],A[2026586:2025078],A[2028095:2026587],tree_1[1350554:1349046],tree_1[1352063:1350555]);
csa_1509 csau_1509_i448(A[2029604:2028096],A[2031113:2029605],A[2032622:2031114],tree_1[1353572:1352064],tree_1[1355081:1353573]);
csa_1509 csau_1509_i449(A[2034131:2032623],A[2035640:2034132],A[2037149:2035641],tree_1[1356590:1355082],tree_1[1358099:1356591]);
csa_1509 csau_1509_i450(A[2038658:2037150],A[2040167:2038659],A[2041676:2040168],tree_1[1359608:1358100],tree_1[1361117:1359609]);
csa_1509 csau_1509_i451(A[2043185:2041677],A[2044694:2043186],A[2046203:2044695],tree_1[1362626:1361118],tree_1[1364135:1362627]);
csa_1509 csau_1509_i452(A[2047712:2046204],A[2049221:2047713],A[2050730:2049222],tree_1[1365644:1364136],tree_1[1367153:1365645]);
csa_1509 csau_1509_i453(A[2052239:2050731],A[2053748:2052240],A[2055257:2053749],tree_1[1368662:1367154],tree_1[1370171:1368663]);
csa_1509 csau_1509_i454(A[2056766:2055258],A[2058275:2056767],A[2059784:2058276],tree_1[1371680:1370172],tree_1[1373189:1371681]);
csa_1509 csau_1509_i455(A[2061293:2059785],A[2062802:2061294],A[2064311:2062803],tree_1[1374698:1373190],tree_1[1376207:1374699]);
csa_1509 csau_1509_i456(A[2065820:2064312],A[2067329:2065821],A[2068838:2067330],tree_1[1377716:1376208],tree_1[1379225:1377717]);
csa_1509 csau_1509_i457(A[2070347:2068839],A[2071856:2070348],A[2073365:2071857],tree_1[1380734:1379226],tree_1[1382243:1380735]);
csa_1509 csau_1509_i458(A[2074874:2073366],A[2076383:2074875],A[2077892:2076384],tree_1[1383752:1382244],tree_1[1385261:1383753]);
csa_1509 csau_1509_i459(A[2079401:2077893],A[2080910:2079402],A[2082419:2080911],tree_1[1386770:1385262],tree_1[1388279:1386771]);
csa_1509 csau_1509_i460(A[2083928:2082420],A[2085437:2083929],A[2086946:2085438],tree_1[1389788:1388280],tree_1[1391297:1389789]);
csa_1509 csau_1509_i461(A[2088455:2086947],A[2089964:2088456],A[2091473:2089965],tree_1[1392806:1391298],tree_1[1394315:1392807]);
csa_1509 csau_1509_i462(A[2092982:2091474],A[2094491:2092983],A[2096000:2094492],tree_1[1395824:1394316],tree_1[1397333:1395825]);
csa_1509 csau_1509_i463(A[2097509:2096001],A[2099018:2097510],A[2100527:2099019],tree_1[1398842:1397334],tree_1[1400351:1398843]);
csa_1509 csau_1509_i464(A[2102036:2100528],A[2103545:2102037],A[2105054:2103546],tree_1[1401860:1400352],tree_1[1403369:1401861]);
csa_1509 csau_1509_i465(A[2106563:2105055],A[2108072:2106564],A[2109581:2108073],tree_1[1404878:1403370],tree_1[1406387:1404879]);
csa_1509 csau_1509_i466(A[2111090:2109582],A[2112599:2111091],A[2114108:2112600],tree_1[1407896:1406388],tree_1[1409405:1407897]);
csa_1509 csau_1509_i467(A[2115617:2114109],A[2117126:2115618],A[2118635:2117127],tree_1[1410914:1409406],tree_1[1412423:1410915]);
csa_1509 csau_1509_i468(A[2120144:2118636],A[2121653:2120145],A[2123162:2121654],tree_1[1413932:1412424],tree_1[1415441:1413933]);
csa_1509 csau_1509_i469(A[2124671:2123163],A[2126180:2124672],A[2127689:2126181],tree_1[1416950:1415442],tree_1[1418459:1416951]);
csa_1509 csau_1509_i470(A[2129198:2127690],A[2130707:2129199],A[2132216:2130708],tree_1[1419968:1418460],tree_1[1421477:1419969]);
csa_1509 csau_1509_i471(A[2133725:2132217],A[2135234:2133726],A[2136743:2135235],tree_1[1422986:1421478],tree_1[1424495:1422987]);
csa_1509 csau_1509_i472(A[2138252:2136744],A[2139761:2138253],A[2141270:2139762],tree_1[1426004:1424496],tree_1[1427513:1426005]);
csa_1509 csau_1509_i473(A[2142779:2141271],A[2144288:2142780],A[2145797:2144289],tree_1[1429022:1427514],tree_1[1430531:1429023]);
csa_1509 csau_1509_i474(A[2147306:2145798],A[2148815:2147307],A[2150324:2148816],tree_1[1432040:1430532],tree_1[1433549:1432041]);
csa_1509 csau_1509_i475(A[2151833:2150325],A[2153342:2151834],A[2154851:2153343],tree_1[1435058:1433550],tree_1[1436567:1435059]);
csa_1509 csau_1509_i476(A[2156360:2154852],A[2157869:2156361],A[2159378:2157870],tree_1[1438076:1436568],tree_1[1439585:1438077]);
csa_1509 csau_1509_i477(A[2160887:2159379],A[2162396:2160888],A[2163905:2162397],tree_1[1441094:1439586],tree_1[1442603:1441095]);
csa_1509 csau_1509_i478(A[2165414:2163906],A[2166923:2165415],A[2168432:2166924],tree_1[1444112:1442604],tree_1[1445621:1444113]);
csa_1509 csau_1509_i479(A[2169941:2168433],A[2171450:2169942],A[2172959:2171451],tree_1[1447130:1445622],tree_1[1448639:1447131]);
csa_1509 csau_1509_i480(A[2174468:2172960],A[2175977:2174469],A[2177486:2175978],tree_1[1450148:1448640],tree_1[1451657:1450149]);
csa_1509 csau_1509_i481(A[2178995:2177487],A[2180504:2178996],A[2182013:2180505],tree_1[1453166:1451658],tree_1[1454675:1453167]);
csa_1509 csau_1509_i482(A[2183522:2182014],A[2185031:2183523],A[2186540:2185032],tree_1[1456184:1454676],tree_1[1457693:1456185]);
csa_1509 csau_1509_i483(A[2188049:2186541],A[2189558:2188050],A[2191067:2189559],tree_1[1459202:1457694],tree_1[1460711:1459203]);
csa_1509 csau_1509_i484(A[2192576:2191068],A[2194085:2192577],A[2195594:2194086],tree_1[1462220:1460712],tree_1[1463729:1462221]);
csa_1509 csau_1509_i485(A[2197103:2195595],A[2198612:2197104],A[2200121:2198613],tree_1[1465238:1463730],tree_1[1466747:1465239]);
csa_1509 csau_1509_i486(A[2201630:2200122],A[2203139:2201631],A[2204648:2203140],tree_1[1468256:1466748],tree_1[1469765:1468257]);
csa_1509 csau_1509_i487(A[2206157:2204649],A[2207666:2206158],A[2209175:2207667],tree_1[1471274:1469766],tree_1[1472783:1471275]);
csa_1509 csau_1509_i488(A[2210684:2209176],A[2212193:2210685],A[2213702:2212194],tree_1[1474292:1472784],tree_1[1475801:1474293]);
csa_1509 csau_1509_i489(A[2215211:2213703],A[2216720:2215212],A[2218229:2216721],tree_1[1477310:1475802],tree_1[1478819:1477311]);
csa_1509 csau_1509_i490(A[2219738:2218230],A[2221247:2219739],A[2222756:2221248],tree_1[1480328:1478820],tree_1[1481837:1480329]);
csa_1509 csau_1509_i491(A[2224265:2222757],A[2225774:2224266],A[2227283:2225775],tree_1[1483346:1481838],tree_1[1484855:1483347]);
csa_1509 csau_1509_i492(A[2228792:2227284],A[2230301:2228793],A[2231810:2230302],tree_1[1486364:1484856],tree_1[1487873:1486365]);
csa_1509 csau_1509_i493(A[2233319:2231811],A[2234828:2233320],A[2236337:2234829],tree_1[1489382:1487874],tree_1[1490891:1489383]);
csa_1509 csau_1509_i494(A[2237846:2236338],A[2239355:2237847],A[2240864:2239356],tree_1[1492400:1490892],tree_1[1493909:1492401]);
csa_1509 csau_1509_i495(A[2242373:2240865],A[2243882:2242374],A[2245391:2243883],tree_1[1495418:1493910],tree_1[1496927:1495419]);
csa_1509 csau_1509_i496(A[2246900:2245392],A[2248409:2246901],A[2249918:2248410],tree_1[1498436:1496928],tree_1[1499945:1498437]);
csa_1509 csau_1509_i497(A[2251427:2249919],A[2252936:2251428],A[2254445:2252937],tree_1[1501454:1499946],tree_1[1502963:1501455]);
csa_1509 csau_1509_i498(A[2255954:2254446],A[2257463:2255955],A[2258972:2257464],tree_1[1504472:1502964],tree_1[1505981:1504473]);
csa_1509 csau_1509_i499(A[2260481:2258973],A[2261990:2260482],A[2263499:2261991],tree_1[1507490:1505982],tree_1[1508999:1507491]);
csa_1509 csau_1509_i500(A[2265008:2263500],A[2266517:2265009],A[2268026:2266518],tree_1[1510508:1509000],tree_1[1512017:1510509]);
csa_1509 csau_1509_i501(A[2269535:2268027],A[2271044:2269536],A[2272553:2271045],tree_1[1513526:1512018],tree_1[1515035:1513527]);
csa_1509 csau_1509_i502(A[2274062:2272554],A[2275571:2274063],A[2277080:2275572],tree_1[1516544:1515036],tree_1[1518053:1516545]);
// layer-2
csa_1509 csau_1509_i503(tree_1[1508:0],tree_1[3017:1509],tree_1[4526:3018],tree_2[1508:0],tree_2[3017:1509]);
csa_1509 csau_1509_i504(tree_1[6035:4527],tree_1[7544:6036],tree_1[9053:7545],tree_2[4526:3018],tree_2[6035:4527]);
csa_1509 csau_1509_i505(tree_1[10562:9054],tree_1[12071:10563],tree_1[13580:12072],tree_2[7544:6036],tree_2[9053:7545]);
csa_1509 csau_1509_i506(tree_1[15089:13581],tree_1[16598:15090],tree_1[18107:16599],tree_2[10562:9054],tree_2[12071:10563]);
csa_1509 csau_1509_i507(tree_1[19616:18108],tree_1[21125:19617],tree_1[22634:21126],tree_2[13580:12072],tree_2[15089:13581]);
csa_1509 csau_1509_i508(tree_1[24143:22635],tree_1[25652:24144],tree_1[27161:25653],tree_2[16598:15090],tree_2[18107:16599]);
csa_1509 csau_1509_i509(tree_1[28670:27162],tree_1[30179:28671],tree_1[31688:30180],tree_2[19616:18108],tree_2[21125:19617]);
csa_1509 csau_1509_i510(tree_1[33197:31689],tree_1[34706:33198],tree_1[36215:34707],tree_2[22634:21126],tree_2[24143:22635]);
csa_1509 csau_1509_i511(tree_1[37724:36216],tree_1[39233:37725],tree_1[40742:39234],tree_2[25652:24144],tree_2[27161:25653]);
csa_1509 csau_1509_i512(tree_1[42251:40743],tree_1[43760:42252],tree_1[45269:43761],tree_2[28670:27162],tree_2[30179:28671]);
csa_1509 csau_1509_i513(tree_1[46778:45270],tree_1[48287:46779],tree_1[49796:48288],tree_2[31688:30180],tree_2[33197:31689]);
csa_1509 csau_1509_i514(tree_1[51305:49797],tree_1[52814:51306],tree_1[54323:52815],tree_2[34706:33198],tree_2[36215:34707]);
csa_1509 csau_1509_i515(tree_1[55832:54324],tree_1[57341:55833],tree_1[58850:57342],tree_2[37724:36216],tree_2[39233:37725]);
csa_1509 csau_1509_i516(tree_1[60359:58851],tree_1[61868:60360],tree_1[63377:61869],tree_2[40742:39234],tree_2[42251:40743]);
csa_1509 csau_1509_i517(tree_1[64886:63378],tree_1[66395:64887],tree_1[67904:66396],tree_2[43760:42252],tree_2[45269:43761]);
csa_1509 csau_1509_i518(tree_1[69413:67905],tree_1[70922:69414],tree_1[72431:70923],tree_2[46778:45270],tree_2[48287:46779]);
csa_1509 csau_1509_i519(tree_1[73940:72432],tree_1[75449:73941],tree_1[76958:75450],tree_2[49796:48288],tree_2[51305:49797]);
csa_1509 csau_1509_i520(tree_1[78467:76959],tree_1[79976:78468],tree_1[81485:79977],tree_2[52814:51306],tree_2[54323:52815]);
csa_1509 csau_1509_i521(tree_1[82994:81486],tree_1[84503:82995],tree_1[86012:84504],tree_2[55832:54324],tree_2[57341:55833]);
csa_1509 csau_1509_i522(tree_1[87521:86013],tree_1[89030:87522],tree_1[90539:89031],tree_2[58850:57342],tree_2[60359:58851]);
csa_1509 csau_1509_i523(tree_1[92048:90540],tree_1[93557:92049],tree_1[95066:93558],tree_2[61868:60360],tree_2[63377:61869]);
csa_1509 csau_1509_i524(tree_1[96575:95067],tree_1[98084:96576],tree_1[99593:98085],tree_2[64886:63378],tree_2[66395:64887]);
csa_1509 csau_1509_i525(tree_1[101102:99594],tree_1[102611:101103],tree_1[104120:102612],tree_2[67904:66396],tree_2[69413:67905]);
csa_1509 csau_1509_i526(tree_1[105629:104121],tree_1[107138:105630],tree_1[108647:107139],tree_2[70922:69414],tree_2[72431:70923]);
csa_1509 csau_1509_i527(tree_1[110156:108648],tree_1[111665:110157],tree_1[113174:111666],tree_2[73940:72432],tree_2[75449:73941]);
csa_1509 csau_1509_i528(tree_1[114683:113175],tree_1[116192:114684],tree_1[117701:116193],tree_2[76958:75450],tree_2[78467:76959]);
csa_1509 csau_1509_i529(tree_1[119210:117702],tree_1[120719:119211],tree_1[122228:120720],tree_2[79976:78468],tree_2[81485:79977]);
csa_1509 csau_1509_i530(tree_1[123737:122229],tree_1[125246:123738],tree_1[126755:125247],tree_2[82994:81486],tree_2[84503:82995]);
csa_1509 csau_1509_i531(tree_1[128264:126756],tree_1[129773:128265],tree_1[131282:129774],tree_2[86012:84504],tree_2[87521:86013]);
csa_1509 csau_1509_i532(tree_1[132791:131283],tree_1[134300:132792],tree_1[135809:134301],tree_2[89030:87522],tree_2[90539:89031]);
csa_1509 csau_1509_i533(tree_1[137318:135810],tree_1[138827:137319],tree_1[140336:138828],tree_2[92048:90540],tree_2[93557:92049]);
csa_1509 csau_1509_i534(tree_1[141845:140337],tree_1[143354:141846],tree_1[144863:143355],tree_2[95066:93558],tree_2[96575:95067]);
csa_1509 csau_1509_i535(tree_1[146372:144864],tree_1[147881:146373],tree_1[149390:147882],tree_2[98084:96576],tree_2[99593:98085]);
csa_1509 csau_1509_i536(tree_1[150899:149391],tree_1[152408:150900],tree_1[153917:152409],tree_2[101102:99594],tree_2[102611:101103]);
csa_1509 csau_1509_i537(tree_1[155426:153918],tree_1[156935:155427],tree_1[158444:156936],tree_2[104120:102612],tree_2[105629:104121]);
csa_1509 csau_1509_i538(tree_1[159953:158445],tree_1[161462:159954],tree_1[162971:161463],tree_2[107138:105630],tree_2[108647:107139]);
csa_1509 csau_1509_i539(tree_1[164480:162972],tree_1[165989:164481],tree_1[167498:165990],tree_2[110156:108648],tree_2[111665:110157]);
csa_1509 csau_1509_i540(tree_1[169007:167499],tree_1[170516:169008],tree_1[172025:170517],tree_2[113174:111666],tree_2[114683:113175]);
csa_1509 csau_1509_i541(tree_1[173534:172026],tree_1[175043:173535],tree_1[176552:175044],tree_2[116192:114684],tree_2[117701:116193]);
csa_1509 csau_1509_i542(tree_1[178061:176553],tree_1[179570:178062],tree_1[181079:179571],tree_2[119210:117702],tree_2[120719:119211]);
csa_1509 csau_1509_i543(tree_1[182588:181080],tree_1[184097:182589],tree_1[185606:184098],tree_2[122228:120720],tree_2[123737:122229]);
csa_1509 csau_1509_i544(tree_1[187115:185607],tree_1[188624:187116],tree_1[190133:188625],tree_2[125246:123738],tree_2[126755:125247]);
csa_1509 csau_1509_i545(tree_1[191642:190134],tree_1[193151:191643],tree_1[194660:193152],tree_2[128264:126756],tree_2[129773:128265]);
csa_1509 csau_1509_i546(tree_1[196169:194661],tree_1[197678:196170],tree_1[199187:197679],tree_2[131282:129774],tree_2[132791:131283]);
csa_1509 csau_1509_i547(tree_1[200696:199188],tree_1[202205:200697],tree_1[203714:202206],tree_2[134300:132792],tree_2[135809:134301]);
csa_1509 csau_1509_i548(tree_1[205223:203715],tree_1[206732:205224],tree_1[208241:206733],tree_2[137318:135810],tree_2[138827:137319]);
csa_1509 csau_1509_i549(tree_1[209750:208242],tree_1[211259:209751],tree_1[212768:211260],tree_2[140336:138828],tree_2[141845:140337]);
csa_1509 csau_1509_i550(tree_1[214277:212769],tree_1[215786:214278],tree_1[217295:215787],tree_2[143354:141846],tree_2[144863:143355]);
csa_1509 csau_1509_i551(tree_1[218804:217296],tree_1[220313:218805],tree_1[221822:220314],tree_2[146372:144864],tree_2[147881:146373]);
csa_1509 csau_1509_i552(tree_1[223331:221823],tree_1[224840:223332],tree_1[226349:224841],tree_2[149390:147882],tree_2[150899:149391]);
csa_1509 csau_1509_i553(tree_1[227858:226350],tree_1[229367:227859],tree_1[230876:229368],tree_2[152408:150900],tree_2[153917:152409]);
csa_1509 csau_1509_i554(tree_1[232385:230877],tree_1[233894:232386],tree_1[235403:233895],tree_2[155426:153918],tree_2[156935:155427]);
csa_1509 csau_1509_i555(tree_1[236912:235404],tree_1[238421:236913],tree_1[239930:238422],tree_2[158444:156936],tree_2[159953:158445]);
csa_1509 csau_1509_i556(tree_1[241439:239931],tree_1[242948:241440],tree_1[244457:242949],tree_2[161462:159954],tree_2[162971:161463]);
csa_1509 csau_1509_i557(tree_1[245966:244458],tree_1[247475:245967],tree_1[248984:247476],tree_2[164480:162972],tree_2[165989:164481]);
csa_1509 csau_1509_i558(tree_1[250493:248985],tree_1[252002:250494],tree_1[253511:252003],tree_2[167498:165990],tree_2[169007:167499]);
csa_1509 csau_1509_i559(tree_1[255020:253512],tree_1[256529:255021],tree_1[258038:256530],tree_2[170516:169008],tree_2[172025:170517]);
csa_1509 csau_1509_i560(tree_1[259547:258039],tree_1[261056:259548],tree_1[262565:261057],tree_2[173534:172026],tree_2[175043:173535]);
csa_1509 csau_1509_i561(tree_1[264074:262566],tree_1[265583:264075],tree_1[267092:265584],tree_2[176552:175044],tree_2[178061:176553]);
csa_1509 csau_1509_i562(tree_1[268601:267093],tree_1[270110:268602],tree_1[271619:270111],tree_2[179570:178062],tree_2[181079:179571]);
csa_1509 csau_1509_i563(tree_1[273128:271620],tree_1[274637:273129],tree_1[276146:274638],tree_2[182588:181080],tree_2[184097:182589]);
csa_1509 csau_1509_i564(tree_1[277655:276147],tree_1[279164:277656],tree_1[280673:279165],tree_2[185606:184098],tree_2[187115:185607]);
csa_1509 csau_1509_i565(tree_1[282182:280674],tree_1[283691:282183],tree_1[285200:283692],tree_2[188624:187116],tree_2[190133:188625]);
csa_1509 csau_1509_i566(tree_1[286709:285201],tree_1[288218:286710],tree_1[289727:288219],tree_2[191642:190134],tree_2[193151:191643]);
csa_1509 csau_1509_i567(tree_1[291236:289728],tree_1[292745:291237],tree_1[294254:292746],tree_2[194660:193152],tree_2[196169:194661]);
csa_1509 csau_1509_i568(tree_1[295763:294255],tree_1[297272:295764],tree_1[298781:297273],tree_2[197678:196170],tree_2[199187:197679]);
csa_1509 csau_1509_i569(tree_1[300290:298782],tree_1[301799:300291],tree_1[303308:301800],tree_2[200696:199188],tree_2[202205:200697]);
csa_1509 csau_1509_i570(tree_1[304817:303309],tree_1[306326:304818],tree_1[307835:306327],tree_2[203714:202206],tree_2[205223:203715]);
csa_1509 csau_1509_i571(tree_1[309344:307836],tree_1[310853:309345],tree_1[312362:310854],tree_2[206732:205224],tree_2[208241:206733]);
csa_1509 csau_1509_i572(tree_1[313871:312363],tree_1[315380:313872],tree_1[316889:315381],tree_2[209750:208242],tree_2[211259:209751]);
csa_1509 csau_1509_i573(tree_1[318398:316890],tree_1[319907:318399],tree_1[321416:319908],tree_2[212768:211260],tree_2[214277:212769]);
csa_1509 csau_1509_i574(tree_1[322925:321417],tree_1[324434:322926],tree_1[325943:324435],tree_2[215786:214278],tree_2[217295:215787]);
csa_1509 csau_1509_i575(tree_1[327452:325944],tree_1[328961:327453],tree_1[330470:328962],tree_2[218804:217296],tree_2[220313:218805]);
csa_1509 csau_1509_i576(tree_1[331979:330471],tree_1[333488:331980],tree_1[334997:333489],tree_2[221822:220314],tree_2[223331:221823]);
csa_1509 csau_1509_i577(tree_1[336506:334998],tree_1[338015:336507],tree_1[339524:338016],tree_2[224840:223332],tree_2[226349:224841]);
csa_1509 csau_1509_i578(tree_1[341033:339525],tree_1[342542:341034],tree_1[344051:342543],tree_2[227858:226350],tree_2[229367:227859]);
csa_1509 csau_1509_i579(tree_1[345560:344052],tree_1[347069:345561],tree_1[348578:347070],tree_2[230876:229368],tree_2[232385:230877]);
csa_1509 csau_1509_i580(tree_1[350087:348579],tree_1[351596:350088],tree_1[353105:351597],tree_2[233894:232386],tree_2[235403:233895]);
csa_1509 csau_1509_i581(tree_1[354614:353106],tree_1[356123:354615],tree_1[357632:356124],tree_2[236912:235404],tree_2[238421:236913]);
csa_1509 csau_1509_i582(tree_1[359141:357633],tree_1[360650:359142],tree_1[362159:360651],tree_2[239930:238422],tree_2[241439:239931]);
csa_1509 csau_1509_i583(tree_1[363668:362160],tree_1[365177:363669],tree_1[366686:365178],tree_2[242948:241440],tree_2[244457:242949]);
csa_1509 csau_1509_i584(tree_1[368195:366687],tree_1[369704:368196],tree_1[371213:369705],tree_2[245966:244458],tree_2[247475:245967]);
csa_1509 csau_1509_i585(tree_1[372722:371214],tree_1[374231:372723],tree_1[375740:374232],tree_2[248984:247476],tree_2[250493:248985]);
csa_1509 csau_1509_i586(tree_1[377249:375741],tree_1[378758:377250],tree_1[380267:378759],tree_2[252002:250494],tree_2[253511:252003]);
csa_1509 csau_1509_i587(tree_1[381776:380268],tree_1[383285:381777],tree_1[384794:383286],tree_2[255020:253512],tree_2[256529:255021]);
csa_1509 csau_1509_i588(tree_1[386303:384795],tree_1[387812:386304],tree_1[389321:387813],tree_2[258038:256530],tree_2[259547:258039]);
csa_1509 csau_1509_i589(tree_1[390830:389322],tree_1[392339:390831],tree_1[393848:392340],tree_2[261056:259548],tree_2[262565:261057]);
csa_1509 csau_1509_i590(tree_1[395357:393849],tree_1[396866:395358],tree_1[398375:396867],tree_2[264074:262566],tree_2[265583:264075]);
csa_1509 csau_1509_i591(tree_1[399884:398376],tree_1[401393:399885],tree_1[402902:401394],tree_2[267092:265584],tree_2[268601:267093]);
csa_1509 csau_1509_i592(tree_1[404411:402903],tree_1[405920:404412],tree_1[407429:405921],tree_2[270110:268602],tree_2[271619:270111]);
csa_1509 csau_1509_i593(tree_1[408938:407430],tree_1[410447:408939],tree_1[411956:410448],tree_2[273128:271620],tree_2[274637:273129]);
csa_1509 csau_1509_i594(tree_1[413465:411957],tree_1[414974:413466],tree_1[416483:414975],tree_2[276146:274638],tree_2[277655:276147]);
csa_1509 csau_1509_i595(tree_1[417992:416484],tree_1[419501:417993],tree_1[421010:419502],tree_2[279164:277656],tree_2[280673:279165]);
csa_1509 csau_1509_i596(tree_1[422519:421011],tree_1[424028:422520],tree_1[425537:424029],tree_2[282182:280674],tree_2[283691:282183]);
csa_1509 csau_1509_i597(tree_1[427046:425538],tree_1[428555:427047],tree_1[430064:428556],tree_2[285200:283692],tree_2[286709:285201]);
csa_1509 csau_1509_i598(tree_1[431573:430065],tree_1[433082:431574],tree_1[434591:433083],tree_2[288218:286710],tree_2[289727:288219]);
csa_1509 csau_1509_i599(tree_1[436100:434592],tree_1[437609:436101],tree_1[439118:437610],tree_2[291236:289728],tree_2[292745:291237]);
csa_1509 csau_1509_i600(tree_1[440627:439119],tree_1[442136:440628],tree_1[443645:442137],tree_2[294254:292746],tree_2[295763:294255]);
csa_1509 csau_1509_i601(tree_1[445154:443646],tree_1[446663:445155],tree_1[448172:446664],tree_2[297272:295764],tree_2[298781:297273]);
csa_1509 csau_1509_i602(tree_1[449681:448173],tree_1[451190:449682],tree_1[452699:451191],tree_2[300290:298782],tree_2[301799:300291]);
csa_1509 csau_1509_i603(tree_1[454208:452700],tree_1[455717:454209],tree_1[457226:455718],tree_2[303308:301800],tree_2[304817:303309]);
csa_1509 csau_1509_i604(tree_1[458735:457227],tree_1[460244:458736],tree_1[461753:460245],tree_2[306326:304818],tree_2[307835:306327]);
csa_1509 csau_1509_i605(tree_1[463262:461754],tree_1[464771:463263],tree_1[466280:464772],tree_2[309344:307836],tree_2[310853:309345]);
csa_1509 csau_1509_i606(tree_1[467789:466281],tree_1[469298:467790],tree_1[470807:469299],tree_2[312362:310854],tree_2[313871:312363]);
csa_1509 csau_1509_i607(tree_1[472316:470808],tree_1[473825:472317],tree_1[475334:473826],tree_2[315380:313872],tree_2[316889:315381]);
csa_1509 csau_1509_i608(tree_1[476843:475335],tree_1[478352:476844],tree_1[479861:478353],tree_2[318398:316890],tree_2[319907:318399]);
csa_1509 csau_1509_i609(tree_1[481370:479862],tree_1[482879:481371],tree_1[484388:482880],tree_2[321416:319908],tree_2[322925:321417]);
csa_1509 csau_1509_i610(tree_1[485897:484389],tree_1[487406:485898],tree_1[488915:487407],tree_2[324434:322926],tree_2[325943:324435]);
csa_1509 csau_1509_i611(tree_1[490424:488916],tree_1[491933:490425],tree_1[493442:491934],tree_2[327452:325944],tree_2[328961:327453]);
csa_1509 csau_1509_i612(tree_1[494951:493443],tree_1[496460:494952],tree_1[497969:496461],tree_2[330470:328962],tree_2[331979:330471]);
csa_1509 csau_1509_i613(tree_1[499478:497970],tree_1[500987:499479],tree_1[502496:500988],tree_2[333488:331980],tree_2[334997:333489]);
csa_1509 csau_1509_i614(tree_1[504005:502497],tree_1[505514:504006],tree_1[507023:505515],tree_2[336506:334998],tree_2[338015:336507]);
csa_1509 csau_1509_i615(tree_1[508532:507024],tree_1[510041:508533],tree_1[511550:510042],tree_2[339524:338016],tree_2[341033:339525]);
csa_1509 csau_1509_i616(tree_1[513059:511551],tree_1[514568:513060],tree_1[516077:514569],tree_2[342542:341034],tree_2[344051:342543]);
csa_1509 csau_1509_i617(tree_1[517586:516078],tree_1[519095:517587],tree_1[520604:519096],tree_2[345560:344052],tree_2[347069:345561]);
csa_1509 csau_1509_i618(tree_1[522113:520605],tree_1[523622:522114],tree_1[525131:523623],tree_2[348578:347070],tree_2[350087:348579]);
csa_1509 csau_1509_i619(tree_1[526640:525132],tree_1[528149:526641],tree_1[529658:528150],tree_2[351596:350088],tree_2[353105:351597]);
csa_1509 csau_1509_i620(tree_1[531167:529659],tree_1[532676:531168],tree_1[534185:532677],tree_2[354614:353106],tree_2[356123:354615]);
csa_1509 csau_1509_i621(tree_1[535694:534186],tree_1[537203:535695],tree_1[538712:537204],tree_2[357632:356124],tree_2[359141:357633]);
csa_1509 csau_1509_i622(tree_1[540221:538713],tree_1[541730:540222],tree_1[543239:541731],tree_2[360650:359142],tree_2[362159:360651]);
csa_1509 csau_1509_i623(tree_1[544748:543240],tree_1[546257:544749],tree_1[547766:546258],tree_2[363668:362160],tree_2[365177:363669]);
csa_1509 csau_1509_i624(tree_1[549275:547767],tree_1[550784:549276],tree_1[552293:550785],tree_2[366686:365178],tree_2[368195:366687]);
csa_1509 csau_1509_i625(tree_1[553802:552294],tree_1[555311:553803],tree_1[556820:555312],tree_2[369704:368196],tree_2[371213:369705]);
csa_1509 csau_1509_i626(tree_1[558329:556821],tree_1[559838:558330],tree_1[561347:559839],tree_2[372722:371214],tree_2[374231:372723]);
csa_1509 csau_1509_i627(tree_1[562856:561348],tree_1[564365:562857],tree_1[565874:564366],tree_2[375740:374232],tree_2[377249:375741]);
csa_1509 csau_1509_i628(tree_1[567383:565875],tree_1[568892:567384],tree_1[570401:568893],tree_2[378758:377250],tree_2[380267:378759]);
csa_1509 csau_1509_i629(tree_1[571910:570402],tree_1[573419:571911],tree_1[574928:573420],tree_2[381776:380268],tree_2[383285:381777]);
csa_1509 csau_1509_i630(tree_1[576437:574929],tree_1[577946:576438],tree_1[579455:577947],tree_2[384794:383286],tree_2[386303:384795]);
csa_1509 csau_1509_i631(tree_1[580964:579456],tree_1[582473:580965],tree_1[583982:582474],tree_2[387812:386304],tree_2[389321:387813]);
csa_1509 csau_1509_i632(tree_1[585491:583983],tree_1[587000:585492],tree_1[588509:587001],tree_2[390830:389322],tree_2[392339:390831]);
csa_1509 csau_1509_i633(tree_1[590018:588510],tree_1[591527:590019],tree_1[593036:591528],tree_2[393848:392340],tree_2[395357:393849]);
csa_1509 csau_1509_i634(tree_1[594545:593037],tree_1[596054:594546],tree_1[597563:596055],tree_2[396866:395358],tree_2[398375:396867]);
csa_1509 csau_1509_i635(tree_1[599072:597564],tree_1[600581:599073],tree_1[602090:600582],tree_2[399884:398376],tree_2[401393:399885]);
csa_1509 csau_1509_i636(tree_1[603599:602091],tree_1[605108:603600],tree_1[606617:605109],tree_2[402902:401394],tree_2[404411:402903]);
csa_1509 csau_1509_i637(tree_1[608126:606618],tree_1[609635:608127],tree_1[611144:609636],tree_2[405920:404412],tree_2[407429:405921]);
csa_1509 csau_1509_i638(tree_1[612653:611145],tree_1[614162:612654],tree_1[615671:614163],tree_2[408938:407430],tree_2[410447:408939]);
csa_1509 csau_1509_i639(tree_1[617180:615672],tree_1[618689:617181],tree_1[620198:618690],tree_2[411956:410448],tree_2[413465:411957]);
csa_1509 csau_1509_i640(tree_1[621707:620199],tree_1[623216:621708],tree_1[624725:623217],tree_2[414974:413466],tree_2[416483:414975]);
csa_1509 csau_1509_i641(tree_1[626234:624726],tree_1[627743:626235],tree_1[629252:627744],tree_2[417992:416484],tree_2[419501:417993]);
csa_1509 csau_1509_i642(tree_1[630761:629253],tree_1[632270:630762],tree_1[633779:632271],tree_2[421010:419502],tree_2[422519:421011]);
csa_1509 csau_1509_i643(tree_1[635288:633780],tree_1[636797:635289],tree_1[638306:636798],tree_2[424028:422520],tree_2[425537:424029]);
csa_1509 csau_1509_i644(tree_1[639815:638307],tree_1[641324:639816],tree_1[642833:641325],tree_2[427046:425538],tree_2[428555:427047]);
csa_1509 csau_1509_i645(tree_1[644342:642834],tree_1[645851:644343],tree_1[647360:645852],tree_2[430064:428556],tree_2[431573:430065]);
csa_1509 csau_1509_i646(tree_1[648869:647361],tree_1[650378:648870],tree_1[651887:650379],tree_2[433082:431574],tree_2[434591:433083]);
csa_1509 csau_1509_i647(tree_1[653396:651888],tree_1[654905:653397],tree_1[656414:654906],tree_2[436100:434592],tree_2[437609:436101]);
csa_1509 csau_1509_i648(tree_1[657923:656415],tree_1[659432:657924],tree_1[660941:659433],tree_2[439118:437610],tree_2[440627:439119]);
csa_1509 csau_1509_i649(tree_1[662450:660942],tree_1[663959:662451],tree_1[665468:663960],tree_2[442136:440628],tree_2[443645:442137]);
csa_1509 csau_1509_i650(tree_1[666977:665469],tree_1[668486:666978],tree_1[669995:668487],tree_2[445154:443646],tree_2[446663:445155]);
csa_1509 csau_1509_i651(tree_1[671504:669996],tree_1[673013:671505],tree_1[674522:673014],tree_2[448172:446664],tree_2[449681:448173]);
csa_1509 csau_1509_i652(tree_1[676031:674523],tree_1[677540:676032],tree_1[679049:677541],tree_2[451190:449682],tree_2[452699:451191]);
csa_1509 csau_1509_i653(tree_1[680558:679050],tree_1[682067:680559],tree_1[683576:682068],tree_2[454208:452700],tree_2[455717:454209]);
csa_1509 csau_1509_i654(tree_1[685085:683577],tree_1[686594:685086],tree_1[688103:686595],tree_2[457226:455718],tree_2[458735:457227]);
csa_1509 csau_1509_i655(tree_1[689612:688104],tree_1[691121:689613],tree_1[692630:691122],tree_2[460244:458736],tree_2[461753:460245]);
csa_1509 csau_1509_i656(tree_1[694139:692631],tree_1[695648:694140],tree_1[697157:695649],tree_2[463262:461754],tree_2[464771:463263]);
csa_1509 csau_1509_i657(tree_1[698666:697158],tree_1[700175:698667],tree_1[701684:700176],tree_2[466280:464772],tree_2[467789:466281]);
csa_1509 csau_1509_i658(tree_1[703193:701685],tree_1[704702:703194],tree_1[706211:704703],tree_2[469298:467790],tree_2[470807:469299]);
csa_1509 csau_1509_i659(tree_1[707720:706212],tree_1[709229:707721],tree_1[710738:709230],tree_2[472316:470808],tree_2[473825:472317]);
csa_1509 csau_1509_i660(tree_1[712247:710739],tree_1[713756:712248],tree_1[715265:713757],tree_2[475334:473826],tree_2[476843:475335]);
csa_1509 csau_1509_i661(tree_1[716774:715266],tree_1[718283:716775],tree_1[719792:718284],tree_2[478352:476844],tree_2[479861:478353]);
csa_1509 csau_1509_i662(tree_1[721301:719793],tree_1[722810:721302],tree_1[724319:722811],tree_2[481370:479862],tree_2[482879:481371]);
csa_1509 csau_1509_i663(tree_1[725828:724320],tree_1[727337:725829],tree_1[728846:727338],tree_2[484388:482880],tree_2[485897:484389]);
csa_1509 csau_1509_i664(tree_1[730355:728847],tree_1[731864:730356],tree_1[733373:731865],tree_2[487406:485898],tree_2[488915:487407]);
csa_1509 csau_1509_i665(tree_1[734882:733374],tree_1[736391:734883],tree_1[737900:736392],tree_2[490424:488916],tree_2[491933:490425]);
csa_1509 csau_1509_i666(tree_1[739409:737901],tree_1[740918:739410],tree_1[742427:740919],tree_2[493442:491934],tree_2[494951:493443]);
csa_1509 csau_1509_i667(tree_1[743936:742428],tree_1[745445:743937],tree_1[746954:745446],tree_2[496460:494952],tree_2[497969:496461]);
csa_1509 csau_1509_i668(tree_1[748463:746955],tree_1[749972:748464],tree_1[751481:749973],tree_2[499478:497970],tree_2[500987:499479]);
csa_1509 csau_1509_i669(tree_1[752990:751482],tree_1[754499:752991],tree_1[756008:754500],tree_2[502496:500988],tree_2[504005:502497]);
csa_1509 csau_1509_i670(tree_1[757517:756009],tree_1[759026:757518],tree_1[760535:759027],tree_2[505514:504006],tree_2[507023:505515]);
csa_1509 csau_1509_i671(tree_1[762044:760536],tree_1[763553:762045],tree_1[765062:763554],tree_2[508532:507024],tree_2[510041:508533]);
csa_1509 csau_1509_i672(tree_1[766571:765063],tree_1[768080:766572],tree_1[769589:768081],tree_2[511550:510042],tree_2[513059:511551]);
csa_1509 csau_1509_i673(tree_1[771098:769590],tree_1[772607:771099],tree_1[774116:772608],tree_2[514568:513060],tree_2[516077:514569]);
csa_1509 csau_1509_i674(tree_1[775625:774117],tree_1[777134:775626],tree_1[778643:777135],tree_2[517586:516078],tree_2[519095:517587]);
csa_1509 csau_1509_i675(tree_1[780152:778644],tree_1[781661:780153],tree_1[783170:781662],tree_2[520604:519096],tree_2[522113:520605]);
csa_1509 csau_1509_i676(tree_1[784679:783171],tree_1[786188:784680],tree_1[787697:786189],tree_2[523622:522114],tree_2[525131:523623]);
csa_1509 csau_1509_i677(tree_1[789206:787698],tree_1[790715:789207],tree_1[792224:790716],tree_2[526640:525132],tree_2[528149:526641]);
csa_1509 csau_1509_i678(tree_1[793733:792225],tree_1[795242:793734],tree_1[796751:795243],tree_2[529658:528150],tree_2[531167:529659]);
csa_1509 csau_1509_i679(tree_1[798260:796752],tree_1[799769:798261],tree_1[801278:799770],tree_2[532676:531168],tree_2[534185:532677]);
csa_1509 csau_1509_i680(tree_1[802787:801279],tree_1[804296:802788],tree_1[805805:804297],tree_2[535694:534186],tree_2[537203:535695]);
csa_1509 csau_1509_i681(tree_1[807314:805806],tree_1[808823:807315],tree_1[810332:808824],tree_2[538712:537204],tree_2[540221:538713]);
csa_1509 csau_1509_i682(tree_1[811841:810333],tree_1[813350:811842],tree_1[814859:813351],tree_2[541730:540222],tree_2[543239:541731]);
csa_1509 csau_1509_i683(tree_1[816368:814860],tree_1[817877:816369],tree_1[819386:817878],tree_2[544748:543240],tree_2[546257:544749]);
csa_1509 csau_1509_i684(tree_1[820895:819387],tree_1[822404:820896],tree_1[823913:822405],tree_2[547766:546258],tree_2[549275:547767]);
csa_1509 csau_1509_i685(tree_1[825422:823914],tree_1[826931:825423],tree_1[828440:826932],tree_2[550784:549276],tree_2[552293:550785]);
csa_1509 csau_1509_i686(tree_1[829949:828441],tree_1[831458:829950],tree_1[832967:831459],tree_2[553802:552294],tree_2[555311:553803]);
csa_1509 csau_1509_i687(tree_1[834476:832968],tree_1[835985:834477],tree_1[837494:835986],tree_2[556820:555312],tree_2[558329:556821]);
csa_1509 csau_1509_i688(tree_1[839003:837495],tree_1[840512:839004],tree_1[842021:840513],tree_2[559838:558330],tree_2[561347:559839]);
csa_1509 csau_1509_i689(tree_1[843530:842022],tree_1[845039:843531],tree_1[846548:845040],tree_2[562856:561348],tree_2[564365:562857]);
csa_1509 csau_1509_i690(tree_1[848057:846549],tree_1[849566:848058],tree_1[851075:849567],tree_2[565874:564366],tree_2[567383:565875]);
csa_1509 csau_1509_i691(tree_1[852584:851076],tree_1[854093:852585],tree_1[855602:854094],tree_2[568892:567384],tree_2[570401:568893]);
csa_1509 csau_1509_i692(tree_1[857111:855603],tree_1[858620:857112],tree_1[860129:858621],tree_2[571910:570402],tree_2[573419:571911]);
csa_1509 csau_1509_i693(tree_1[861638:860130],tree_1[863147:861639],tree_1[864656:863148],tree_2[574928:573420],tree_2[576437:574929]);
csa_1509 csau_1509_i694(tree_1[866165:864657],tree_1[867674:866166],tree_1[869183:867675],tree_2[577946:576438],tree_2[579455:577947]);
csa_1509 csau_1509_i695(tree_1[870692:869184],tree_1[872201:870693],tree_1[873710:872202],tree_2[580964:579456],tree_2[582473:580965]);
csa_1509 csau_1509_i696(tree_1[875219:873711],tree_1[876728:875220],tree_1[878237:876729],tree_2[583982:582474],tree_2[585491:583983]);
csa_1509 csau_1509_i697(tree_1[879746:878238],tree_1[881255:879747],tree_1[882764:881256],tree_2[587000:585492],tree_2[588509:587001]);
csa_1509 csau_1509_i698(tree_1[884273:882765],tree_1[885782:884274],tree_1[887291:885783],tree_2[590018:588510],tree_2[591527:590019]);
csa_1509 csau_1509_i699(tree_1[888800:887292],tree_1[890309:888801],tree_1[891818:890310],tree_2[593036:591528],tree_2[594545:593037]);
csa_1509 csau_1509_i700(tree_1[893327:891819],tree_1[894836:893328],tree_1[896345:894837],tree_2[596054:594546],tree_2[597563:596055]);
csa_1509 csau_1509_i701(tree_1[897854:896346],tree_1[899363:897855],tree_1[900872:899364],tree_2[599072:597564],tree_2[600581:599073]);
csa_1509 csau_1509_i702(tree_1[902381:900873],tree_1[903890:902382],tree_1[905399:903891],tree_2[602090:600582],tree_2[603599:602091]);
csa_1509 csau_1509_i703(tree_1[906908:905400],tree_1[908417:906909],tree_1[909926:908418],tree_2[605108:603600],tree_2[606617:605109]);
csa_1509 csau_1509_i704(tree_1[911435:909927],tree_1[912944:911436],tree_1[914453:912945],tree_2[608126:606618],tree_2[609635:608127]);
csa_1509 csau_1509_i705(tree_1[915962:914454],tree_1[917471:915963],tree_1[918980:917472],tree_2[611144:609636],tree_2[612653:611145]);
csa_1509 csau_1509_i706(tree_1[920489:918981],tree_1[921998:920490],tree_1[923507:921999],tree_2[614162:612654],tree_2[615671:614163]);
csa_1509 csau_1509_i707(tree_1[925016:923508],tree_1[926525:925017],tree_1[928034:926526],tree_2[617180:615672],tree_2[618689:617181]);
csa_1509 csau_1509_i708(tree_1[929543:928035],tree_1[931052:929544],tree_1[932561:931053],tree_2[620198:618690],tree_2[621707:620199]);
csa_1509 csau_1509_i709(tree_1[934070:932562],tree_1[935579:934071],tree_1[937088:935580],tree_2[623216:621708],tree_2[624725:623217]);
csa_1509 csau_1509_i710(tree_1[938597:937089],tree_1[940106:938598],tree_1[941615:940107],tree_2[626234:624726],tree_2[627743:626235]);
csa_1509 csau_1509_i711(tree_1[943124:941616],tree_1[944633:943125],tree_1[946142:944634],tree_2[629252:627744],tree_2[630761:629253]);
csa_1509 csau_1509_i712(tree_1[947651:946143],tree_1[949160:947652],tree_1[950669:949161],tree_2[632270:630762],tree_2[633779:632271]);
csa_1509 csau_1509_i713(tree_1[952178:950670],tree_1[953687:952179],tree_1[955196:953688],tree_2[635288:633780],tree_2[636797:635289]);
csa_1509 csau_1509_i714(tree_1[956705:955197],tree_1[958214:956706],tree_1[959723:958215],tree_2[638306:636798],tree_2[639815:638307]);
csa_1509 csau_1509_i715(tree_1[961232:959724],tree_1[962741:961233],tree_1[964250:962742],tree_2[641324:639816],tree_2[642833:641325]);
csa_1509 csau_1509_i716(tree_1[965759:964251],tree_1[967268:965760],tree_1[968777:967269],tree_2[644342:642834],tree_2[645851:644343]);
csa_1509 csau_1509_i717(tree_1[970286:968778],tree_1[971795:970287],tree_1[973304:971796],tree_2[647360:645852],tree_2[648869:647361]);
csa_1509 csau_1509_i718(tree_1[974813:973305],tree_1[976322:974814],tree_1[977831:976323],tree_2[650378:648870],tree_2[651887:650379]);
csa_1509 csau_1509_i719(tree_1[979340:977832],tree_1[980849:979341],tree_1[982358:980850],tree_2[653396:651888],tree_2[654905:653397]);
csa_1509 csau_1509_i720(tree_1[983867:982359],tree_1[985376:983868],tree_1[986885:985377],tree_2[656414:654906],tree_2[657923:656415]);
csa_1509 csau_1509_i721(tree_1[988394:986886],tree_1[989903:988395],tree_1[991412:989904],tree_2[659432:657924],tree_2[660941:659433]);
csa_1509 csau_1509_i722(tree_1[992921:991413],tree_1[994430:992922],tree_1[995939:994431],tree_2[662450:660942],tree_2[663959:662451]);
csa_1509 csau_1509_i723(tree_1[997448:995940],tree_1[998957:997449],tree_1[1000466:998958],tree_2[665468:663960],tree_2[666977:665469]);
csa_1509 csau_1509_i724(tree_1[1001975:1000467],tree_1[1003484:1001976],tree_1[1004993:1003485],tree_2[668486:666978],tree_2[669995:668487]);
csa_1509 csau_1509_i725(tree_1[1006502:1004994],tree_1[1008011:1006503],tree_1[1009520:1008012],tree_2[671504:669996],tree_2[673013:671505]);
csa_1509 csau_1509_i726(tree_1[1011029:1009521],tree_1[1012538:1011030],tree_1[1014047:1012539],tree_2[674522:673014],tree_2[676031:674523]);
csa_1509 csau_1509_i727(tree_1[1015556:1014048],tree_1[1017065:1015557],tree_1[1018574:1017066],tree_2[677540:676032],tree_2[679049:677541]);
csa_1509 csau_1509_i728(tree_1[1020083:1018575],tree_1[1021592:1020084],tree_1[1023101:1021593],tree_2[680558:679050],tree_2[682067:680559]);
csa_1509 csau_1509_i729(tree_1[1024610:1023102],tree_1[1026119:1024611],tree_1[1027628:1026120],tree_2[683576:682068],tree_2[685085:683577]);
csa_1509 csau_1509_i730(tree_1[1029137:1027629],tree_1[1030646:1029138],tree_1[1032155:1030647],tree_2[686594:685086],tree_2[688103:686595]);
csa_1509 csau_1509_i731(tree_1[1033664:1032156],tree_1[1035173:1033665],tree_1[1036682:1035174],tree_2[689612:688104],tree_2[691121:689613]);
csa_1509 csau_1509_i732(tree_1[1038191:1036683],tree_1[1039700:1038192],tree_1[1041209:1039701],tree_2[692630:691122],tree_2[694139:692631]);
csa_1509 csau_1509_i733(tree_1[1042718:1041210],tree_1[1044227:1042719],tree_1[1045736:1044228],tree_2[695648:694140],tree_2[697157:695649]);
csa_1509 csau_1509_i734(tree_1[1047245:1045737],tree_1[1048754:1047246],tree_1[1050263:1048755],tree_2[698666:697158],tree_2[700175:698667]);
csa_1509 csau_1509_i735(tree_1[1051772:1050264],tree_1[1053281:1051773],tree_1[1054790:1053282],tree_2[701684:700176],tree_2[703193:701685]);
csa_1509 csau_1509_i736(tree_1[1056299:1054791],tree_1[1057808:1056300],tree_1[1059317:1057809],tree_2[704702:703194],tree_2[706211:704703]);
csa_1509 csau_1509_i737(tree_1[1060826:1059318],tree_1[1062335:1060827],tree_1[1063844:1062336],tree_2[707720:706212],tree_2[709229:707721]);
csa_1509 csau_1509_i738(tree_1[1065353:1063845],tree_1[1066862:1065354],tree_1[1068371:1066863],tree_2[710738:709230],tree_2[712247:710739]);
csa_1509 csau_1509_i739(tree_1[1069880:1068372],tree_1[1071389:1069881],tree_1[1072898:1071390],tree_2[713756:712248],tree_2[715265:713757]);
csa_1509 csau_1509_i740(tree_1[1074407:1072899],tree_1[1075916:1074408],tree_1[1077425:1075917],tree_2[716774:715266],tree_2[718283:716775]);
csa_1509 csau_1509_i741(tree_1[1078934:1077426],tree_1[1080443:1078935],tree_1[1081952:1080444],tree_2[719792:718284],tree_2[721301:719793]);
csa_1509 csau_1509_i742(tree_1[1083461:1081953],tree_1[1084970:1083462],tree_1[1086479:1084971],tree_2[722810:721302],tree_2[724319:722811]);
csa_1509 csau_1509_i743(tree_1[1087988:1086480],tree_1[1089497:1087989],tree_1[1091006:1089498],tree_2[725828:724320],tree_2[727337:725829]);
csa_1509 csau_1509_i744(tree_1[1092515:1091007],tree_1[1094024:1092516],tree_1[1095533:1094025],tree_2[728846:727338],tree_2[730355:728847]);
csa_1509 csau_1509_i745(tree_1[1097042:1095534],tree_1[1098551:1097043],tree_1[1100060:1098552],tree_2[731864:730356],tree_2[733373:731865]);
csa_1509 csau_1509_i746(tree_1[1101569:1100061],tree_1[1103078:1101570],tree_1[1104587:1103079],tree_2[734882:733374],tree_2[736391:734883]);
csa_1509 csau_1509_i747(tree_1[1106096:1104588],tree_1[1107605:1106097],tree_1[1109114:1107606],tree_2[737900:736392],tree_2[739409:737901]);
csa_1509 csau_1509_i748(tree_1[1110623:1109115],tree_1[1112132:1110624],tree_1[1113641:1112133],tree_2[740918:739410],tree_2[742427:740919]);
csa_1509 csau_1509_i749(tree_1[1115150:1113642],tree_1[1116659:1115151],tree_1[1118168:1116660],tree_2[743936:742428],tree_2[745445:743937]);
csa_1509 csau_1509_i750(tree_1[1119677:1118169],tree_1[1121186:1119678],tree_1[1122695:1121187],tree_2[746954:745446],tree_2[748463:746955]);
csa_1509 csau_1509_i751(tree_1[1124204:1122696],tree_1[1125713:1124205],tree_1[1127222:1125714],tree_2[749972:748464],tree_2[751481:749973]);
csa_1509 csau_1509_i752(tree_1[1128731:1127223],tree_1[1130240:1128732],tree_1[1131749:1130241],tree_2[752990:751482],tree_2[754499:752991]);
csa_1509 csau_1509_i753(tree_1[1133258:1131750],tree_1[1134767:1133259],tree_1[1136276:1134768],tree_2[756008:754500],tree_2[757517:756009]);
csa_1509 csau_1509_i754(tree_1[1137785:1136277],tree_1[1139294:1137786],tree_1[1140803:1139295],tree_2[759026:757518],tree_2[760535:759027]);
csa_1509 csau_1509_i755(tree_1[1142312:1140804],tree_1[1143821:1142313],tree_1[1145330:1143822],tree_2[762044:760536],tree_2[763553:762045]);
csa_1509 csau_1509_i756(tree_1[1146839:1145331],tree_1[1148348:1146840],tree_1[1149857:1148349],tree_2[765062:763554],tree_2[766571:765063]);
csa_1509 csau_1509_i757(tree_1[1151366:1149858],tree_1[1152875:1151367],tree_1[1154384:1152876],tree_2[768080:766572],tree_2[769589:768081]);
csa_1509 csau_1509_i758(tree_1[1155893:1154385],tree_1[1157402:1155894],tree_1[1158911:1157403],tree_2[771098:769590],tree_2[772607:771099]);
csa_1509 csau_1509_i759(tree_1[1160420:1158912],tree_1[1161929:1160421],tree_1[1163438:1161930],tree_2[774116:772608],tree_2[775625:774117]);
csa_1509 csau_1509_i760(tree_1[1164947:1163439],tree_1[1166456:1164948],tree_1[1167965:1166457],tree_2[777134:775626],tree_2[778643:777135]);
csa_1509 csau_1509_i761(tree_1[1169474:1167966],tree_1[1170983:1169475],tree_1[1172492:1170984],tree_2[780152:778644],tree_2[781661:780153]);
csa_1509 csau_1509_i762(tree_1[1174001:1172493],tree_1[1175510:1174002],tree_1[1177019:1175511],tree_2[783170:781662],tree_2[784679:783171]);
csa_1509 csau_1509_i763(tree_1[1178528:1177020],tree_1[1180037:1178529],tree_1[1181546:1180038],tree_2[786188:784680],tree_2[787697:786189]);
csa_1509 csau_1509_i764(tree_1[1183055:1181547],tree_1[1184564:1183056],tree_1[1186073:1184565],tree_2[789206:787698],tree_2[790715:789207]);
csa_1509 csau_1509_i765(tree_1[1187582:1186074],tree_1[1189091:1187583],tree_1[1190600:1189092],tree_2[792224:790716],tree_2[793733:792225]);
csa_1509 csau_1509_i766(tree_1[1192109:1190601],tree_1[1193618:1192110],tree_1[1195127:1193619],tree_2[795242:793734],tree_2[796751:795243]);
csa_1509 csau_1509_i767(tree_1[1196636:1195128],tree_1[1198145:1196637],tree_1[1199654:1198146],tree_2[798260:796752],tree_2[799769:798261]);
csa_1509 csau_1509_i768(tree_1[1201163:1199655],tree_1[1202672:1201164],tree_1[1204181:1202673],tree_2[801278:799770],tree_2[802787:801279]);
csa_1509 csau_1509_i769(tree_1[1205690:1204182],tree_1[1207199:1205691],tree_1[1208708:1207200],tree_2[804296:802788],tree_2[805805:804297]);
csa_1509 csau_1509_i770(tree_1[1210217:1208709],tree_1[1211726:1210218],tree_1[1213235:1211727],tree_2[807314:805806],tree_2[808823:807315]);
csa_1509 csau_1509_i771(tree_1[1214744:1213236],tree_1[1216253:1214745],tree_1[1217762:1216254],tree_2[810332:808824],tree_2[811841:810333]);
csa_1509 csau_1509_i772(tree_1[1219271:1217763],tree_1[1220780:1219272],tree_1[1222289:1220781],tree_2[813350:811842],tree_2[814859:813351]);
csa_1509 csau_1509_i773(tree_1[1223798:1222290],tree_1[1225307:1223799],tree_1[1226816:1225308],tree_2[816368:814860],tree_2[817877:816369]);
csa_1509 csau_1509_i774(tree_1[1228325:1226817],tree_1[1229834:1228326],tree_1[1231343:1229835],tree_2[819386:817878],tree_2[820895:819387]);
csa_1509 csau_1509_i775(tree_1[1232852:1231344],tree_1[1234361:1232853],tree_1[1235870:1234362],tree_2[822404:820896],tree_2[823913:822405]);
csa_1509 csau_1509_i776(tree_1[1237379:1235871],tree_1[1238888:1237380],tree_1[1240397:1238889],tree_2[825422:823914],tree_2[826931:825423]);
csa_1509 csau_1509_i777(tree_1[1241906:1240398],tree_1[1243415:1241907],tree_1[1244924:1243416],tree_2[828440:826932],tree_2[829949:828441]);
csa_1509 csau_1509_i778(tree_1[1246433:1244925],tree_1[1247942:1246434],tree_1[1249451:1247943],tree_2[831458:829950],tree_2[832967:831459]);
csa_1509 csau_1509_i779(tree_1[1250960:1249452],tree_1[1252469:1250961],tree_1[1253978:1252470],tree_2[834476:832968],tree_2[835985:834477]);
csa_1509 csau_1509_i780(tree_1[1255487:1253979],tree_1[1256996:1255488],tree_1[1258505:1256997],tree_2[837494:835986],tree_2[839003:837495]);
csa_1509 csau_1509_i781(tree_1[1260014:1258506],tree_1[1261523:1260015],tree_1[1263032:1261524],tree_2[840512:839004],tree_2[842021:840513]);
csa_1509 csau_1509_i782(tree_1[1264541:1263033],tree_1[1266050:1264542],tree_1[1267559:1266051],tree_2[843530:842022],tree_2[845039:843531]);
csa_1509 csau_1509_i783(tree_1[1269068:1267560],tree_1[1270577:1269069],tree_1[1272086:1270578],tree_2[846548:845040],tree_2[848057:846549]);
csa_1509 csau_1509_i784(tree_1[1273595:1272087],tree_1[1275104:1273596],tree_1[1276613:1275105],tree_2[849566:848058],tree_2[851075:849567]);
csa_1509 csau_1509_i785(tree_1[1278122:1276614],tree_1[1279631:1278123],tree_1[1281140:1279632],tree_2[852584:851076],tree_2[854093:852585]);
csa_1509 csau_1509_i786(tree_1[1282649:1281141],tree_1[1284158:1282650],tree_1[1285667:1284159],tree_2[855602:854094],tree_2[857111:855603]);
csa_1509 csau_1509_i787(tree_1[1287176:1285668],tree_1[1288685:1287177],tree_1[1290194:1288686],tree_2[858620:857112],tree_2[860129:858621]);
csa_1509 csau_1509_i788(tree_1[1291703:1290195],tree_1[1293212:1291704],tree_1[1294721:1293213],tree_2[861638:860130],tree_2[863147:861639]);
csa_1509 csau_1509_i789(tree_1[1296230:1294722],tree_1[1297739:1296231],tree_1[1299248:1297740],tree_2[864656:863148],tree_2[866165:864657]);
csa_1509 csau_1509_i790(tree_1[1300757:1299249],tree_1[1302266:1300758],tree_1[1303775:1302267],tree_2[867674:866166],tree_2[869183:867675]);
csa_1509 csau_1509_i791(tree_1[1305284:1303776],tree_1[1306793:1305285],tree_1[1308302:1306794],tree_2[870692:869184],tree_2[872201:870693]);
csa_1509 csau_1509_i792(tree_1[1309811:1308303],tree_1[1311320:1309812],tree_1[1312829:1311321],tree_2[873710:872202],tree_2[875219:873711]);
csa_1509 csau_1509_i793(tree_1[1314338:1312830],tree_1[1315847:1314339],tree_1[1317356:1315848],tree_2[876728:875220],tree_2[878237:876729]);
csa_1509 csau_1509_i794(tree_1[1318865:1317357],tree_1[1320374:1318866],tree_1[1321883:1320375],tree_2[879746:878238],tree_2[881255:879747]);
csa_1509 csau_1509_i795(tree_1[1323392:1321884],tree_1[1324901:1323393],tree_1[1326410:1324902],tree_2[882764:881256],tree_2[884273:882765]);
csa_1509 csau_1509_i796(tree_1[1327919:1326411],tree_1[1329428:1327920],tree_1[1330937:1329429],tree_2[885782:884274],tree_2[887291:885783]);
csa_1509 csau_1509_i797(tree_1[1332446:1330938],tree_1[1333955:1332447],tree_1[1335464:1333956],tree_2[888800:887292],tree_2[890309:888801]);
csa_1509 csau_1509_i798(tree_1[1336973:1335465],tree_1[1338482:1336974],tree_1[1339991:1338483],tree_2[891818:890310],tree_2[893327:891819]);
csa_1509 csau_1509_i799(tree_1[1341500:1339992],tree_1[1343009:1341501],tree_1[1344518:1343010],tree_2[894836:893328],tree_2[896345:894837]);
csa_1509 csau_1509_i800(tree_1[1346027:1344519],tree_1[1347536:1346028],tree_1[1349045:1347537],tree_2[897854:896346],tree_2[899363:897855]);
csa_1509 csau_1509_i801(tree_1[1350554:1349046],tree_1[1352063:1350555],tree_1[1353572:1352064],tree_2[900872:899364],tree_2[902381:900873]);
csa_1509 csau_1509_i802(tree_1[1355081:1353573],tree_1[1356590:1355082],tree_1[1358099:1356591],tree_2[903890:902382],tree_2[905399:903891]);
csa_1509 csau_1509_i803(tree_1[1359608:1358100],tree_1[1361117:1359609],tree_1[1362626:1361118],tree_2[906908:905400],tree_2[908417:906909]);
csa_1509 csau_1509_i804(tree_1[1364135:1362627],tree_1[1365644:1364136],tree_1[1367153:1365645],tree_2[909926:908418],tree_2[911435:909927]);
csa_1509 csau_1509_i805(tree_1[1368662:1367154],tree_1[1370171:1368663],tree_1[1371680:1370172],tree_2[912944:911436],tree_2[914453:912945]);
csa_1509 csau_1509_i806(tree_1[1373189:1371681],tree_1[1374698:1373190],tree_1[1376207:1374699],tree_2[915962:914454],tree_2[917471:915963]);
csa_1509 csau_1509_i807(tree_1[1377716:1376208],tree_1[1379225:1377717],tree_1[1380734:1379226],tree_2[918980:917472],tree_2[920489:918981]);
csa_1509 csau_1509_i808(tree_1[1382243:1380735],tree_1[1383752:1382244],tree_1[1385261:1383753],tree_2[921998:920490],tree_2[923507:921999]);
csa_1509 csau_1509_i809(tree_1[1386770:1385262],tree_1[1388279:1386771],tree_1[1389788:1388280],tree_2[925016:923508],tree_2[926525:925017]);
csa_1509 csau_1509_i810(tree_1[1391297:1389789],tree_1[1392806:1391298],tree_1[1394315:1392807],tree_2[928034:926526],tree_2[929543:928035]);
csa_1509 csau_1509_i811(tree_1[1395824:1394316],tree_1[1397333:1395825],tree_1[1398842:1397334],tree_2[931052:929544],tree_2[932561:931053]);
csa_1509 csau_1509_i812(tree_1[1400351:1398843],tree_1[1401860:1400352],tree_1[1403369:1401861],tree_2[934070:932562],tree_2[935579:934071]);
csa_1509 csau_1509_i813(tree_1[1404878:1403370],tree_1[1406387:1404879],tree_1[1407896:1406388],tree_2[937088:935580],tree_2[938597:937089]);
csa_1509 csau_1509_i814(tree_1[1409405:1407897],tree_1[1410914:1409406],tree_1[1412423:1410915],tree_2[940106:938598],tree_2[941615:940107]);
csa_1509 csau_1509_i815(tree_1[1413932:1412424],tree_1[1415441:1413933],tree_1[1416950:1415442],tree_2[943124:941616],tree_2[944633:943125]);
csa_1509 csau_1509_i816(tree_1[1418459:1416951],tree_1[1419968:1418460],tree_1[1421477:1419969],tree_2[946142:944634],tree_2[947651:946143]);
csa_1509 csau_1509_i817(tree_1[1422986:1421478],tree_1[1424495:1422987],tree_1[1426004:1424496],tree_2[949160:947652],tree_2[950669:949161]);
csa_1509 csau_1509_i818(tree_1[1427513:1426005],tree_1[1429022:1427514],tree_1[1430531:1429023],tree_2[952178:950670],tree_2[953687:952179]);
csa_1509 csau_1509_i819(tree_1[1432040:1430532],tree_1[1433549:1432041],tree_1[1435058:1433550],tree_2[955196:953688],tree_2[956705:955197]);
csa_1509 csau_1509_i820(tree_1[1436567:1435059],tree_1[1438076:1436568],tree_1[1439585:1438077],tree_2[958214:956706],tree_2[959723:958215]);
csa_1509 csau_1509_i821(tree_1[1441094:1439586],tree_1[1442603:1441095],tree_1[1444112:1442604],tree_2[961232:959724],tree_2[962741:961233]);
csa_1509 csau_1509_i822(tree_1[1445621:1444113],tree_1[1447130:1445622],tree_1[1448639:1447131],tree_2[964250:962742],tree_2[965759:964251]);
csa_1509 csau_1509_i823(tree_1[1450148:1448640],tree_1[1451657:1450149],tree_1[1453166:1451658],tree_2[967268:965760],tree_2[968777:967269]);
csa_1509 csau_1509_i824(tree_1[1454675:1453167],tree_1[1456184:1454676],tree_1[1457693:1456185],tree_2[970286:968778],tree_2[971795:970287]);
csa_1509 csau_1509_i825(tree_1[1459202:1457694],tree_1[1460711:1459203],tree_1[1462220:1460712],tree_2[973304:971796],tree_2[974813:973305]);
csa_1509 csau_1509_i826(tree_1[1463729:1462221],tree_1[1465238:1463730],tree_1[1466747:1465239],tree_2[976322:974814],tree_2[977831:976323]);
csa_1509 csau_1509_i827(tree_1[1468256:1466748],tree_1[1469765:1468257],tree_1[1471274:1469766],tree_2[979340:977832],tree_2[980849:979341]);
csa_1509 csau_1509_i828(tree_1[1472783:1471275],tree_1[1474292:1472784],tree_1[1475801:1474293],tree_2[982358:980850],tree_2[983867:982359]);
csa_1509 csau_1509_i829(tree_1[1477310:1475802],tree_1[1478819:1477311],tree_1[1480328:1478820],tree_2[985376:983868],tree_2[986885:985377]);
csa_1509 csau_1509_i830(tree_1[1481837:1480329],tree_1[1483346:1481838],tree_1[1484855:1483347],tree_2[988394:986886],tree_2[989903:988395]);
csa_1509 csau_1509_i831(tree_1[1486364:1484856],tree_1[1487873:1486365],tree_1[1489382:1487874],tree_2[991412:989904],tree_2[992921:991413]);
csa_1509 csau_1509_i832(tree_1[1490891:1489383],tree_1[1492400:1490892],tree_1[1493909:1492401],tree_2[994430:992922],tree_2[995939:994431]);
csa_1509 csau_1509_i833(tree_1[1495418:1493910],tree_1[1496927:1495419],tree_1[1498436:1496928],tree_2[997448:995940],tree_2[998957:997449]);
csa_1509 csau_1509_i834(tree_1[1499945:1498437],tree_1[1501454:1499946],tree_1[1502963:1501455],tree_2[1000466:998958],tree_2[1001975:1000467]);
csa_1509 csau_1509_i835(tree_1[1504472:1502964],tree_1[1505981:1504473],tree_1[1507490:1505982],tree_2[1003484:1001976],tree_2[1004993:1003485]);
csa_1509 csau_1509_i836(tree_1[1508999:1507491],tree_1[1510508:1509000],tree_1[1512017:1510509],tree_2[1006502:1004994],tree_2[1008011:1006503]);
csa_1509 csau_1509_i837(tree_1[1513526:1512018],tree_1[1515035:1513527],tree_1[1516544:1515036],tree_2[1009520:1008012],tree_2[1011029:1009521]);
assign tree_2[1012538:1011030] = tree_1[1518053:1516545];
// layer-3
csa_1509 csau_1509_i838(tree_2[1508:0],tree_2[3017:1509],tree_2[4526:3018],tree_3[1508:0],tree_3[3017:1509]);
csa_1509 csau_1509_i839(tree_2[6035:4527],tree_2[7544:6036],tree_2[9053:7545],tree_3[4526:3018],tree_3[6035:4527]);
csa_1509 csau_1509_i840(tree_2[10562:9054],tree_2[12071:10563],tree_2[13580:12072],tree_3[7544:6036],tree_3[9053:7545]);
csa_1509 csau_1509_i841(tree_2[15089:13581],tree_2[16598:15090],tree_2[18107:16599],tree_3[10562:9054],tree_3[12071:10563]);
csa_1509 csau_1509_i842(tree_2[19616:18108],tree_2[21125:19617],tree_2[22634:21126],tree_3[13580:12072],tree_3[15089:13581]);
csa_1509 csau_1509_i843(tree_2[24143:22635],tree_2[25652:24144],tree_2[27161:25653],tree_3[16598:15090],tree_3[18107:16599]);
csa_1509 csau_1509_i844(tree_2[28670:27162],tree_2[30179:28671],tree_2[31688:30180],tree_3[19616:18108],tree_3[21125:19617]);
csa_1509 csau_1509_i845(tree_2[33197:31689],tree_2[34706:33198],tree_2[36215:34707],tree_3[22634:21126],tree_3[24143:22635]);
csa_1509 csau_1509_i846(tree_2[37724:36216],tree_2[39233:37725],tree_2[40742:39234],tree_3[25652:24144],tree_3[27161:25653]);
csa_1509 csau_1509_i847(tree_2[42251:40743],tree_2[43760:42252],tree_2[45269:43761],tree_3[28670:27162],tree_3[30179:28671]);
csa_1509 csau_1509_i848(tree_2[46778:45270],tree_2[48287:46779],tree_2[49796:48288],tree_3[31688:30180],tree_3[33197:31689]);
csa_1509 csau_1509_i849(tree_2[51305:49797],tree_2[52814:51306],tree_2[54323:52815],tree_3[34706:33198],tree_3[36215:34707]);
csa_1509 csau_1509_i850(tree_2[55832:54324],tree_2[57341:55833],tree_2[58850:57342],tree_3[37724:36216],tree_3[39233:37725]);
csa_1509 csau_1509_i851(tree_2[60359:58851],tree_2[61868:60360],tree_2[63377:61869],tree_3[40742:39234],tree_3[42251:40743]);
csa_1509 csau_1509_i852(tree_2[64886:63378],tree_2[66395:64887],tree_2[67904:66396],tree_3[43760:42252],tree_3[45269:43761]);
csa_1509 csau_1509_i853(tree_2[69413:67905],tree_2[70922:69414],tree_2[72431:70923],tree_3[46778:45270],tree_3[48287:46779]);
csa_1509 csau_1509_i854(tree_2[73940:72432],tree_2[75449:73941],tree_2[76958:75450],tree_3[49796:48288],tree_3[51305:49797]);
csa_1509 csau_1509_i855(tree_2[78467:76959],tree_2[79976:78468],tree_2[81485:79977],tree_3[52814:51306],tree_3[54323:52815]);
csa_1509 csau_1509_i856(tree_2[82994:81486],tree_2[84503:82995],tree_2[86012:84504],tree_3[55832:54324],tree_3[57341:55833]);
csa_1509 csau_1509_i857(tree_2[87521:86013],tree_2[89030:87522],tree_2[90539:89031],tree_3[58850:57342],tree_3[60359:58851]);
csa_1509 csau_1509_i858(tree_2[92048:90540],tree_2[93557:92049],tree_2[95066:93558],tree_3[61868:60360],tree_3[63377:61869]);
csa_1509 csau_1509_i859(tree_2[96575:95067],tree_2[98084:96576],tree_2[99593:98085],tree_3[64886:63378],tree_3[66395:64887]);
csa_1509 csau_1509_i860(tree_2[101102:99594],tree_2[102611:101103],tree_2[104120:102612],tree_3[67904:66396],tree_3[69413:67905]);
csa_1509 csau_1509_i861(tree_2[105629:104121],tree_2[107138:105630],tree_2[108647:107139],tree_3[70922:69414],tree_3[72431:70923]);
csa_1509 csau_1509_i862(tree_2[110156:108648],tree_2[111665:110157],tree_2[113174:111666],tree_3[73940:72432],tree_3[75449:73941]);
csa_1509 csau_1509_i863(tree_2[114683:113175],tree_2[116192:114684],tree_2[117701:116193],tree_3[76958:75450],tree_3[78467:76959]);
csa_1509 csau_1509_i864(tree_2[119210:117702],tree_2[120719:119211],tree_2[122228:120720],tree_3[79976:78468],tree_3[81485:79977]);
csa_1509 csau_1509_i865(tree_2[123737:122229],tree_2[125246:123738],tree_2[126755:125247],tree_3[82994:81486],tree_3[84503:82995]);
csa_1509 csau_1509_i866(tree_2[128264:126756],tree_2[129773:128265],tree_2[131282:129774],tree_3[86012:84504],tree_3[87521:86013]);
csa_1509 csau_1509_i867(tree_2[132791:131283],tree_2[134300:132792],tree_2[135809:134301],tree_3[89030:87522],tree_3[90539:89031]);
csa_1509 csau_1509_i868(tree_2[137318:135810],tree_2[138827:137319],tree_2[140336:138828],tree_3[92048:90540],tree_3[93557:92049]);
csa_1509 csau_1509_i869(tree_2[141845:140337],tree_2[143354:141846],tree_2[144863:143355],tree_3[95066:93558],tree_3[96575:95067]);
csa_1509 csau_1509_i870(tree_2[146372:144864],tree_2[147881:146373],tree_2[149390:147882],tree_3[98084:96576],tree_3[99593:98085]);
csa_1509 csau_1509_i871(tree_2[150899:149391],tree_2[152408:150900],tree_2[153917:152409],tree_3[101102:99594],tree_3[102611:101103]);
csa_1509 csau_1509_i872(tree_2[155426:153918],tree_2[156935:155427],tree_2[158444:156936],tree_3[104120:102612],tree_3[105629:104121]);
csa_1509 csau_1509_i873(tree_2[159953:158445],tree_2[161462:159954],tree_2[162971:161463],tree_3[107138:105630],tree_3[108647:107139]);
csa_1509 csau_1509_i874(tree_2[164480:162972],tree_2[165989:164481],tree_2[167498:165990],tree_3[110156:108648],tree_3[111665:110157]);
csa_1509 csau_1509_i875(tree_2[169007:167499],tree_2[170516:169008],tree_2[172025:170517],tree_3[113174:111666],tree_3[114683:113175]);
csa_1509 csau_1509_i876(tree_2[173534:172026],tree_2[175043:173535],tree_2[176552:175044],tree_3[116192:114684],tree_3[117701:116193]);
csa_1509 csau_1509_i877(tree_2[178061:176553],tree_2[179570:178062],tree_2[181079:179571],tree_3[119210:117702],tree_3[120719:119211]);
csa_1509 csau_1509_i878(tree_2[182588:181080],tree_2[184097:182589],tree_2[185606:184098],tree_3[122228:120720],tree_3[123737:122229]);
csa_1509 csau_1509_i879(tree_2[187115:185607],tree_2[188624:187116],tree_2[190133:188625],tree_3[125246:123738],tree_3[126755:125247]);
csa_1509 csau_1509_i880(tree_2[191642:190134],tree_2[193151:191643],tree_2[194660:193152],tree_3[128264:126756],tree_3[129773:128265]);
csa_1509 csau_1509_i881(tree_2[196169:194661],tree_2[197678:196170],tree_2[199187:197679],tree_3[131282:129774],tree_3[132791:131283]);
csa_1509 csau_1509_i882(tree_2[200696:199188],tree_2[202205:200697],tree_2[203714:202206],tree_3[134300:132792],tree_3[135809:134301]);
csa_1509 csau_1509_i883(tree_2[205223:203715],tree_2[206732:205224],tree_2[208241:206733],tree_3[137318:135810],tree_3[138827:137319]);
csa_1509 csau_1509_i884(tree_2[209750:208242],tree_2[211259:209751],tree_2[212768:211260],tree_3[140336:138828],tree_3[141845:140337]);
csa_1509 csau_1509_i885(tree_2[214277:212769],tree_2[215786:214278],tree_2[217295:215787],tree_3[143354:141846],tree_3[144863:143355]);
csa_1509 csau_1509_i886(tree_2[218804:217296],tree_2[220313:218805],tree_2[221822:220314],tree_3[146372:144864],tree_3[147881:146373]);
csa_1509 csau_1509_i887(tree_2[223331:221823],tree_2[224840:223332],tree_2[226349:224841],tree_3[149390:147882],tree_3[150899:149391]);
csa_1509 csau_1509_i888(tree_2[227858:226350],tree_2[229367:227859],tree_2[230876:229368],tree_3[152408:150900],tree_3[153917:152409]);
csa_1509 csau_1509_i889(tree_2[232385:230877],tree_2[233894:232386],tree_2[235403:233895],tree_3[155426:153918],tree_3[156935:155427]);
csa_1509 csau_1509_i890(tree_2[236912:235404],tree_2[238421:236913],tree_2[239930:238422],tree_3[158444:156936],tree_3[159953:158445]);
csa_1509 csau_1509_i891(tree_2[241439:239931],tree_2[242948:241440],tree_2[244457:242949],tree_3[161462:159954],tree_3[162971:161463]);
csa_1509 csau_1509_i892(tree_2[245966:244458],tree_2[247475:245967],tree_2[248984:247476],tree_3[164480:162972],tree_3[165989:164481]);
csa_1509 csau_1509_i893(tree_2[250493:248985],tree_2[252002:250494],tree_2[253511:252003],tree_3[167498:165990],tree_3[169007:167499]);
csa_1509 csau_1509_i894(tree_2[255020:253512],tree_2[256529:255021],tree_2[258038:256530],tree_3[170516:169008],tree_3[172025:170517]);
csa_1509 csau_1509_i895(tree_2[259547:258039],tree_2[261056:259548],tree_2[262565:261057],tree_3[173534:172026],tree_3[175043:173535]);
csa_1509 csau_1509_i896(tree_2[264074:262566],tree_2[265583:264075],tree_2[267092:265584],tree_3[176552:175044],tree_3[178061:176553]);
csa_1509 csau_1509_i897(tree_2[268601:267093],tree_2[270110:268602],tree_2[271619:270111],tree_3[179570:178062],tree_3[181079:179571]);
csa_1509 csau_1509_i898(tree_2[273128:271620],tree_2[274637:273129],tree_2[276146:274638],tree_3[182588:181080],tree_3[184097:182589]);
csa_1509 csau_1509_i899(tree_2[277655:276147],tree_2[279164:277656],tree_2[280673:279165],tree_3[185606:184098],tree_3[187115:185607]);
csa_1509 csau_1509_i900(tree_2[282182:280674],tree_2[283691:282183],tree_2[285200:283692],tree_3[188624:187116],tree_3[190133:188625]);
csa_1509 csau_1509_i901(tree_2[286709:285201],tree_2[288218:286710],tree_2[289727:288219],tree_3[191642:190134],tree_3[193151:191643]);
csa_1509 csau_1509_i902(tree_2[291236:289728],tree_2[292745:291237],tree_2[294254:292746],tree_3[194660:193152],tree_3[196169:194661]);
csa_1509 csau_1509_i903(tree_2[295763:294255],tree_2[297272:295764],tree_2[298781:297273],tree_3[197678:196170],tree_3[199187:197679]);
csa_1509 csau_1509_i904(tree_2[300290:298782],tree_2[301799:300291],tree_2[303308:301800],tree_3[200696:199188],tree_3[202205:200697]);
csa_1509 csau_1509_i905(tree_2[304817:303309],tree_2[306326:304818],tree_2[307835:306327],tree_3[203714:202206],tree_3[205223:203715]);
csa_1509 csau_1509_i906(tree_2[309344:307836],tree_2[310853:309345],tree_2[312362:310854],tree_3[206732:205224],tree_3[208241:206733]);
csa_1509 csau_1509_i907(tree_2[313871:312363],tree_2[315380:313872],tree_2[316889:315381],tree_3[209750:208242],tree_3[211259:209751]);
csa_1509 csau_1509_i908(tree_2[318398:316890],tree_2[319907:318399],tree_2[321416:319908],tree_3[212768:211260],tree_3[214277:212769]);
csa_1509 csau_1509_i909(tree_2[322925:321417],tree_2[324434:322926],tree_2[325943:324435],tree_3[215786:214278],tree_3[217295:215787]);
csa_1509 csau_1509_i910(tree_2[327452:325944],tree_2[328961:327453],tree_2[330470:328962],tree_3[218804:217296],tree_3[220313:218805]);
csa_1509 csau_1509_i911(tree_2[331979:330471],tree_2[333488:331980],tree_2[334997:333489],tree_3[221822:220314],tree_3[223331:221823]);
csa_1509 csau_1509_i912(tree_2[336506:334998],tree_2[338015:336507],tree_2[339524:338016],tree_3[224840:223332],tree_3[226349:224841]);
csa_1509 csau_1509_i913(tree_2[341033:339525],tree_2[342542:341034],tree_2[344051:342543],tree_3[227858:226350],tree_3[229367:227859]);
csa_1509 csau_1509_i914(tree_2[345560:344052],tree_2[347069:345561],tree_2[348578:347070],tree_3[230876:229368],tree_3[232385:230877]);
csa_1509 csau_1509_i915(tree_2[350087:348579],tree_2[351596:350088],tree_2[353105:351597],tree_3[233894:232386],tree_3[235403:233895]);
csa_1509 csau_1509_i916(tree_2[354614:353106],tree_2[356123:354615],tree_2[357632:356124],tree_3[236912:235404],tree_3[238421:236913]);
csa_1509 csau_1509_i917(tree_2[359141:357633],tree_2[360650:359142],tree_2[362159:360651],tree_3[239930:238422],tree_3[241439:239931]);
csa_1509 csau_1509_i918(tree_2[363668:362160],tree_2[365177:363669],tree_2[366686:365178],tree_3[242948:241440],tree_3[244457:242949]);
csa_1509 csau_1509_i919(tree_2[368195:366687],tree_2[369704:368196],tree_2[371213:369705],tree_3[245966:244458],tree_3[247475:245967]);
csa_1509 csau_1509_i920(tree_2[372722:371214],tree_2[374231:372723],tree_2[375740:374232],tree_3[248984:247476],tree_3[250493:248985]);
csa_1509 csau_1509_i921(tree_2[377249:375741],tree_2[378758:377250],tree_2[380267:378759],tree_3[252002:250494],tree_3[253511:252003]);
csa_1509 csau_1509_i922(tree_2[381776:380268],tree_2[383285:381777],tree_2[384794:383286],tree_3[255020:253512],tree_3[256529:255021]);
csa_1509 csau_1509_i923(tree_2[386303:384795],tree_2[387812:386304],tree_2[389321:387813],tree_3[258038:256530],tree_3[259547:258039]);
csa_1509 csau_1509_i924(tree_2[390830:389322],tree_2[392339:390831],tree_2[393848:392340],tree_3[261056:259548],tree_3[262565:261057]);
csa_1509 csau_1509_i925(tree_2[395357:393849],tree_2[396866:395358],tree_2[398375:396867],tree_3[264074:262566],tree_3[265583:264075]);
csa_1509 csau_1509_i926(tree_2[399884:398376],tree_2[401393:399885],tree_2[402902:401394],tree_3[267092:265584],tree_3[268601:267093]);
csa_1509 csau_1509_i927(tree_2[404411:402903],tree_2[405920:404412],tree_2[407429:405921],tree_3[270110:268602],tree_3[271619:270111]);
csa_1509 csau_1509_i928(tree_2[408938:407430],tree_2[410447:408939],tree_2[411956:410448],tree_3[273128:271620],tree_3[274637:273129]);
csa_1509 csau_1509_i929(tree_2[413465:411957],tree_2[414974:413466],tree_2[416483:414975],tree_3[276146:274638],tree_3[277655:276147]);
csa_1509 csau_1509_i930(tree_2[417992:416484],tree_2[419501:417993],tree_2[421010:419502],tree_3[279164:277656],tree_3[280673:279165]);
csa_1509 csau_1509_i931(tree_2[422519:421011],tree_2[424028:422520],tree_2[425537:424029],tree_3[282182:280674],tree_3[283691:282183]);
csa_1509 csau_1509_i932(tree_2[427046:425538],tree_2[428555:427047],tree_2[430064:428556],tree_3[285200:283692],tree_3[286709:285201]);
csa_1509 csau_1509_i933(tree_2[431573:430065],tree_2[433082:431574],tree_2[434591:433083],tree_3[288218:286710],tree_3[289727:288219]);
csa_1509 csau_1509_i934(tree_2[436100:434592],tree_2[437609:436101],tree_2[439118:437610],tree_3[291236:289728],tree_3[292745:291237]);
csa_1509 csau_1509_i935(tree_2[440627:439119],tree_2[442136:440628],tree_2[443645:442137],tree_3[294254:292746],tree_3[295763:294255]);
csa_1509 csau_1509_i936(tree_2[445154:443646],tree_2[446663:445155],tree_2[448172:446664],tree_3[297272:295764],tree_3[298781:297273]);
csa_1509 csau_1509_i937(tree_2[449681:448173],tree_2[451190:449682],tree_2[452699:451191],tree_3[300290:298782],tree_3[301799:300291]);
csa_1509 csau_1509_i938(tree_2[454208:452700],tree_2[455717:454209],tree_2[457226:455718],tree_3[303308:301800],tree_3[304817:303309]);
csa_1509 csau_1509_i939(tree_2[458735:457227],tree_2[460244:458736],tree_2[461753:460245],tree_3[306326:304818],tree_3[307835:306327]);
csa_1509 csau_1509_i940(tree_2[463262:461754],tree_2[464771:463263],tree_2[466280:464772],tree_3[309344:307836],tree_3[310853:309345]);
csa_1509 csau_1509_i941(tree_2[467789:466281],tree_2[469298:467790],tree_2[470807:469299],tree_3[312362:310854],tree_3[313871:312363]);
csa_1509 csau_1509_i942(tree_2[472316:470808],tree_2[473825:472317],tree_2[475334:473826],tree_3[315380:313872],tree_3[316889:315381]);
csa_1509 csau_1509_i943(tree_2[476843:475335],tree_2[478352:476844],tree_2[479861:478353],tree_3[318398:316890],tree_3[319907:318399]);
csa_1509 csau_1509_i944(tree_2[481370:479862],tree_2[482879:481371],tree_2[484388:482880],tree_3[321416:319908],tree_3[322925:321417]);
csa_1509 csau_1509_i945(tree_2[485897:484389],tree_2[487406:485898],tree_2[488915:487407],tree_3[324434:322926],tree_3[325943:324435]);
csa_1509 csau_1509_i946(tree_2[490424:488916],tree_2[491933:490425],tree_2[493442:491934],tree_3[327452:325944],tree_3[328961:327453]);
csa_1509 csau_1509_i947(tree_2[494951:493443],tree_2[496460:494952],tree_2[497969:496461],tree_3[330470:328962],tree_3[331979:330471]);
csa_1509 csau_1509_i948(tree_2[499478:497970],tree_2[500987:499479],tree_2[502496:500988],tree_3[333488:331980],tree_3[334997:333489]);
csa_1509 csau_1509_i949(tree_2[504005:502497],tree_2[505514:504006],tree_2[507023:505515],tree_3[336506:334998],tree_3[338015:336507]);
csa_1509 csau_1509_i950(tree_2[508532:507024],tree_2[510041:508533],tree_2[511550:510042],tree_3[339524:338016],tree_3[341033:339525]);
csa_1509 csau_1509_i951(tree_2[513059:511551],tree_2[514568:513060],tree_2[516077:514569],tree_3[342542:341034],tree_3[344051:342543]);
csa_1509 csau_1509_i952(tree_2[517586:516078],tree_2[519095:517587],tree_2[520604:519096],tree_3[345560:344052],tree_3[347069:345561]);
csa_1509 csau_1509_i953(tree_2[522113:520605],tree_2[523622:522114],tree_2[525131:523623],tree_3[348578:347070],tree_3[350087:348579]);
csa_1509 csau_1509_i954(tree_2[526640:525132],tree_2[528149:526641],tree_2[529658:528150],tree_3[351596:350088],tree_3[353105:351597]);
csa_1509 csau_1509_i955(tree_2[531167:529659],tree_2[532676:531168],tree_2[534185:532677],tree_3[354614:353106],tree_3[356123:354615]);
csa_1509 csau_1509_i956(tree_2[535694:534186],tree_2[537203:535695],tree_2[538712:537204],tree_3[357632:356124],tree_3[359141:357633]);
csa_1509 csau_1509_i957(tree_2[540221:538713],tree_2[541730:540222],tree_2[543239:541731],tree_3[360650:359142],tree_3[362159:360651]);
csa_1509 csau_1509_i958(tree_2[544748:543240],tree_2[546257:544749],tree_2[547766:546258],tree_3[363668:362160],tree_3[365177:363669]);
csa_1509 csau_1509_i959(tree_2[549275:547767],tree_2[550784:549276],tree_2[552293:550785],tree_3[366686:365178],tree_3[368195:366687]);
csa_1509 csau_1509_i960(tree_2[553802:552294],tree_2[555311:553803],tree_2[556820:555312],tree_3[369704:368196],tree_3[371213:369705]);
csa_1509 csau_1509_i961(tree_2[558329:556821],tree_2[559838:558330],tree_2[561347:559839],tree_3[372722:371214],tree_3[374231:372723]);
csa_1509 csau_1509_i962(tree_2[562856:561348],tree_2[564365:562857],tree_2[565874:564366],tree_3[375740:374232],tree_3[377249:375741]);
csa_1509 csau_1509_i963(tree_2[567383:565875],tree_2[568892:567384],tree_2[570401:568893],tree_3[378758:377250],tree_3[380267:378759]);
csa_1509 csau_1509_i964(tree_2[571910:570402],tree_2[573419:571911],tree_2[574928:573420],tree_3[381776:380268],tree_3[383285:381777]);
csa_1509 csau_1509_i965(tree_2[576437:574929],tree_2[577946:576438],tree_2[579455:577947],tree_3[384794:383286],tree_3[386303:384795]);
csa_1509 csau_1509_i966(tree_2[580964:579456],tree_2[582473:580965],tree_2[583982:582474],tree_3[387812:386304],tree_3[389321:387813]);
csa_1509 csau_1509_i967(tree_2[585491:583983],tree_2[587000:585492],tree_2[588509:587001],tree_3[390830:389322],tree_3[392339:390831]);
csa_1509 csau_1509_i968(tree_2[590018:588510],tree_2[591527:590019],tree_2[593036:591528],tree_3[393848:392340],tree_3[395357:393849]);
csa_1509 csau_1509_i969(tree_2[594545:593037],tree_2[596054:594546],tree_2[597563:596055],tree_3[396866:395358],tree_3[398375:396867]);
csa_1509 csau_1509_i970(tree_2[599072:597564],tree_2[600581:599073],tree_2[602090:600582],tree_3[399884:398376],tree_3[401393:399885]);
csa_1509 csau_1509_i971(tree_2[603599:602091],tree_2[605108:603600],tree_2[606617:605109],tree_3[402902:401394],tree_3[404411:402903]);
csa_1509 csau_1509_i972(tree_2[608126:606618],tree_2[609635:608127],tree_2[611144:609636],tree_3[405920:404412],tree_3[407429:405921]);
csa_1509 csau_1509_i973(tree_2[612653:611145],tree_2[614162:612654],tree_2[615671:614163],tree_3[408938:407430],tree_3[410447:408939]);
csa_1509 csau_1509_i974(tree_2[617180:615672],tree_2[618689:617181],tree_2[620198:618690],tree_3[411956:410448],tree_3[413465:411957]);
csa_1509 csau_1509_i975(tree_2[621707:620199],tree_2[623216:621708],tree_2[624725:623217],tree_3[414974:413466],tree_3[416483:414975]);
csa_1509 csau_1509_i976(tree_2[626234:624726],tree_2[627743:626235],tree_2[629252:627744],tree_3[417992:416484],tree_3[419501:417993]);
csa_1509 csau_1509_i977(tree_2[630761:629253],tree_2[632270:630762],tree_2[633779:632271],tree_3[421010:419502],tree_3[422519:421011]);
csa_1509 csau_1509_i978(tree_2[635288:633780],tree_2[636797:635289],tree_2[638306:636798],tree_3[424028:422520],tree_3[425537:424029]);
csa_1509 csau_1509_i979(tree_2[639815:638307],tree_2[641324:639816],tree_2[642833:641325],tree_3[427046:425538],tree_3[428555:427047]);
csa_1509 csau_1509_i980(tree_2[644342:642834],tree_2[645851:644343],tree_2[647360:645852],tree_3[430064:428556],tree_3[431573:430065]);
csa_1509 csau_1509_i981(tree_2[648869:647361],tree_2[650378:648870],tree_2[651887:650379],tree_3[433082:431574],tree_3[434591:433083]);
csa_1509 csau_1509_i982(tree_2[653396:651888],tree_2[654905:653397],tree_2[656414:654906],tree_3[436100:434592],tree_3[437609:436101]);
csa_1509 csau_1509_i983(tree_2[657923:656415],tree_2[659432:657924],tree_2[660941:659433],tree_3[439118:437610],tree_3[440627:439119]);
csa_1509 csau_1509_i984(tree_2[662450:660942],tree_2[663959:662451],tree_2[665468:663960],tree_3[442136:440628],tree_3[443645:442137]);
csa_1509 csau_1509_i985(tree_2[666977:665469],tree_2[668486:666978],tree_2[669995:668487],tree_3[445154:443646],tree_3[446663:445155]);
csa_1509 csau_1509_i986(tree_2[671504:669996],tree_2[673013:671505],tree_2[674522:673014],tree_3[448172:446664],tree_3[449681:448173]);
csa_1509 csau_1509_i987(tree_2[676031:674523],tree_2[677540:676032],tree_2[679049:677541],tree_3[451190:449682],tree_3[452699:451191]);
csa_1509 csau_1509_i988(tree_2[680558:679050],tree_2[682067:680559],tree_2[683576:682068],tree_3[454208:452700],tree_3[455717:454209]);
csa_1509 csau_1509_i989(tree_2[685085:683577],tree_2[686594:685086],tree_2[688103:686595],tree_3[457226:455718],tree_3[458735:457227]);
csa_1509 csau_1509_i990(tree_2[689612:688104],tree_2[691121:689613],tree_2[692630:691122],tree_3[460244:458736],tree_3[461753:460245]);
csa_1509 csau_1509_i991(tree_2[694139:692631],tree_2[695648:694140],tree_2[697157:695649],tree_3[463262:461754],tree_3[464771:463263]);
csa_1509 csau_1509_i992(tree_2[698666:697158],tree_2[700175:698667],tree_2[701684:700176],tree_3[466280:464772],tree_3[467789:466281]);
csa_1509 csau_1509_i993(tree_2[703193:701685],tree_2[704702:703194],tree_2[706211:704703],tree_3[469298:467790],tree_3[470807:469299]);
csa_1509 csau_1509_i994(tree_2[707720:706212],tree_2[709229:707721],tree_2[710738:709230],tree_3[472316:470808],tree_3[473825:472317]);
csa_1509 csau_1509_i995(tree_2[712247:710739],tree_2[713756:712248],tree_2[715265:713757],tree_3[475334:473826],tree_3[476843:475335]);
csa_1509 csau_1509_i996(tree_2[716774:715266],tree_2[718283:716775],tree_2[719792:718284],tree_3[478352:476844],tree_3[479861:478353]);
csa_1509 csau_1509_i997(tree_2[721301:719793],tree_2[722810:721302],tree_2[724319:722811],tree_3[481370:479862],tree_3[482879:481371]);
csa_1509 csau_1509_i998(tree_2[725828:724320],tree_2[727337:725829],tree_2[728846:727338],tree_3[484388:482880],tree_3[485897:484389]);
csa_1509 csau_1509_i999(tree_2[730355:728847],tree_2[731864:730356],tree_2[733373:731865],tree_3[487406:485898],tree_3[488915:487407]);
csa_1509 csau_1509_i1000(tree_2[734882:733374],tree_2[736391:734883],tree_2[737900:736392],tree_3[490424:488916],tree_3[491933:490425]);
csa_1509 csau_1509_i1001(tree_2[739409:737901],tree_2[740918:739410],tree_2[742427:740919],tree_3[493442:491934],tree_3[494951:493443]);
csa_1509 csau_1509_i1002(tree_2[743936:742428],tree_2[745445:743937],tree_2[746954:745446],tree_3[496460:494952],tree_3[497969:496461]);
csa_1509 csau_1509_i1003(tree_2[748463:746955],tree_2[749972:748464],tree_2[751481:749973],tree_3[499478:497970],tree_3[500987:499479]);
csa_1509 csau_1509_i1004(tree_2[752990:751482],tree_2[754499:752991],tree_2[756008:754500],tree_3[502496:500988],tree_3[504005:502497]);
csa_1509 csau_1509_i1005(tree_2[757517:756009],tree_2[759026:757518],tree_2[760535:759027],tree_3[505514:504006],tree_3[507023:505515]);
csa_1509 csau_1509_i1006(tree_2[762044:760536],tree_2[763553:762045],tree_2[765062:763554],tree_3[508532:507024],tree_3[510041:508533]);
csa_1509 csau_1509_i1007(tree_2[766571:765063],tree_2[768080:766572],tree_2[769589:768081],tree_3[511550:510042],tree_3[513059:511551]);
csa_1509 csau_1509_i1008(tree_2[771098:769590],tree_2[772607:771099],tree_2[774116:772608],tree_3[514568:513060],tree_3[516077:514569]);
csa_1509 csau_1509_i1009(tree_2[775625:774117],tree_2[777134:775626],tree_2[778643:777135],tree_3[517586:516078],tree_3[519095:517587]);
csa_1509 csau_1509_i1010(tree_2[780152:778644],tree_2[781661:780153],tree_2[783170:781662],tree_3[520604:519096],tree_3[522113:520605]);
csa_1509 csau_1509_i1011(tree_2[784679:783171],tree_2[786188:784680],tree_2[787697:786189],tree_3[523622:522114],tree_3[525131:523623]);
csa_1509 csau_1509_i1012(tree_2[789206:787698],tree_2[790715:789207],tree_2[792224:790716],tree_3[526640:525132],tree_3[528149:526641]);
csa_1509 csau_1509_i1013(tree_2[793733:792225],tree_2[795242:793734],tree_2[796751:795243],tree_3[529658:528150],tree_3[531167:529659]);
csa_1509 csau_1509_i1014(tree_2[798260:796752],tree_2[799769:798261],tree_2[801278:799770],tree_3[532676:531168],tree_3[534185:532677]);
csa_1509 csau_1509_i1015(tree_2[802787:801279],tree_2[804296:802788],tree_2[805805:804297],tree_3[535694:534186],tree_3[537203:535695]);
csa_1509 csau_1509_i1016(tree_2[807314:805806],tree_2[808823:807315],tree_2[810332:808824],tree_3[538712:537204],tree_3[540221:538713]);
csa_1509 csau_1509_i1017(tree_2[811841:810333],tree_2[813350:811842],tree_2[814859:813351],tree_3[541730:540222],tree_3[543239:541731]);
csa_1509 csau_1509_i1018(tree_2[816368:814860],tree_2[817877:816369],tree_2[819386:817878],tree_3[544748:543240],tree_3[546257:544749]);
csa_1509 csau_1509_i1019(tree_2[820895:819387],tree_2[822404:820896],tree_2[823913:822405],tree_3[547766:546258],tree_3[549275:547767]);
csa_1509 csau_1509_i1020(tree_2[825422:823914],tree_2[826931:825423],tree_2[828440:826932],tree_3[550784:549276],tree_3[552293:550785]);
csa_1509 csau_1509_i1021(tree_2[829949:828441],tree_2[831458:829950],tree_2[832967:831459],tree_3[553802:552294],tree_3[555311:553803]);
csa_1509 csau_1509_i1022(tree_2[834476:832968],tree_2[835985:834477],tree_2[837494:835986],tree_3[556820:555312],tree_3[558329:556821]);
csa_1509 csau_1509_i1023(tree_2[839003:837495],tree_2[840512:839004],tree_2[842021:840513],tree_3[559838:558330],tree_3[561347:559839]);
csa_1509 csau_1509_i1024(tree_2[843530:842022],tree_2[845039:843531],tree_2[846548:845040],tree_3[562856:561348],tree_3[564365:562857]);
csa_1509 csau_1509_i1025(tree_2[848057:846549],tree_2[849566:848058],tree_2[851075:849567],tree_3[565874:564366],tree_3[567383:565875]);
csa_1509 csau_1509_i1026(tree_2[852584:851076],tree_2[854093:852585],tree_2[855602:854094],tree_3[568892:567384],tree_3[570401:568893]);
csa_1509 csau_1509_i1027(tree_2[857111:855603],tree_2[858620:857112],tree_2[860129:858621],tree_3[571910:570402],tree_3[573419:571911]);
csa_1509 csau_1509_i1028(tree_2[861638:860130],tree_2[863147:861639],tree_2[864656:863148],tree_3[574928:573420],tree_3[576437:574929]);
csa_1509 csau_1509_i1029(tree_2[866165:864657],tree_2[867674:866166],tree_2[869183:867675],tree_3[577946:576438],tree_3[579455:577947]);
csa_1509 csau_1509_i1030(tree_2[870692:869184],tree_2[872201:870693],tree_2[873710:872202],tree_3[580964:579456],tree_3[582473:580965]);
csa_1509 csau_1509_i1031(tree_2[875219:873711],tree_2[876728:875220],tree_2[878237:876729],tree_3[583982:582474],tree_3[585491:583983]);
csa_1509 csau_1509_i1032(tree_2[879746:878238],tree_2[881255:879747],tree_2[882764:881256],tree_3[587000:585492],tree_3[588509:587001]);
csa_1509 csau_1509_i1033(tree_2[884273:882765],tree_2[885782:884274],tree_2[887291:885783],tree_3[590018:588510],tree_3[591527:590019]);
csa_1509 csau_1509_i1034(tree_2[888800:887292],tree_2[890309:888801],tree_2[891818:890310],tree_3[593036:591528],tree_3[594545:593037]);
csa_1509 csau_1509_i1035(tree_2[893327:891819],tree_2[894836:893328],tree_2[896345:894837],tree_3[596054:594546],tree_3[597563:596055]);
csa_1509 csau_1509_i1036(tree_2[897854:896346],tree_2[899363:897855],tree_2[900872:899364],tree_3[599072:597564],tree_3[600581:599073]);
csa_1509 csau_1509_i1037(tree_2[902381:900873],tree_2[903890:902382],tree_2[905399:903891],tree_3[602090:600582],tree_3[603599:602091]);
csa_1509 csau_1509_i1038(tree_2[906908:905400],tree_2[908417:906909],tree_2[909926:908418],tree_3[605108:603600],tree_3[606617:605109]);
csa_1509 csau_1509_i1039(tree_2[911435:909927],tree_2[912944:911436],tree_2[914453:912945],tree_3[608126:606618],tree_3[609635:608127]);
csa_1509 csau_1509_i1040(tree_2[915962:914454],tree_2[917471:915963],tree_2[918980:917472],tree_3[611144:609636],tree_3[612653:611145]);
csa_1509 csau_1509_i1041(tree_2[920489:918981],tree_2[921998:920490],tree_2[923507:921999],tree_3[614162:612654],tree_3[615671:614163]);
csa_1509 csau_1509_i1042(tree_2[925016:923508],tree_2[926525:925017],tree_2[928034:926526],tree_3[617180:615672],tree_3[618689:617181]);
csa_1509 csau_1509_i1043(tree_2[929543:928035],tree_2[931052:929544],tree_2[932561:931053],tree_3[620198:618690],tree_3[621707:620199]);
csa_1509 csau_1509_i1044(tree_2[934070:932562],tree_2[935579:934071],tree_2[937088:935580],tree_3[623216:621708],tree_3[624725:623217]);
csa_1509 csau_1509_i1045(tree_2[938597:937089],tree_2[940106:938598],tree_2[941615:940107],tree_3[626234:624726],tree_3[627743:626235]);
csa_1509 csau_1509_i1046(tree_2[943124:941616],tree_2[944633:943125],tree_2[946142:944634],tree_3[629252:627744],tree_3[630761:629253]);
csa_1509 csau_1509_i1047(tree_2[947651:946143],tree_2[949160:947652],tree_2[950669:949161],tree_3[632270:630762],tree_3[633779:632271]);
csa_1509 csau_1509_i1048(tree_2[952178:950670],tree_2[953687:952179],tree_2[955196:953688],tree_3[635288:633780],tree_3[636797:635289]);
csa_1509 csau_1509_i1049(tree_2[956705:955197],tree_2[958214:956706],tree_2[959723:958215],tree_3[638306:636798],tree_3[639815:638307]);
csa_1509 csau_1509_i1050(tree_2[961232:959724],tree_2[962741:961233],tree_2[964250:962742],tree_3[641324:639816],tree_3[642833:641325]);
csa_1509 csau_1509_i1051(tree_2[965759:964251],tree_2[967268:965760],tree_2[968777:967269],tree_3[644342:642834],tree_3[645851:644343]);
csa_1509 csau_1509_i1052(tree_2[970286:968778],tree_2[971795:970287],tree_2[973304:971796],tree_3[647360:645852],tree_3[648869:647361]);
csa_1509 csau_1509_i1053(tree_2[974813:973305],tree_2[976322:974814],tree_2[977831:976323],tree_3[650378:648870],tree_3[651887:650379]);
csa_1509 csau_1509_i1054(tree_2[979340:977832],tree_2[980849:979341],tree_2[982358:980850],tree_3[653396:651888],tree_3[654905:653397]);
csa_1509 csau_1509_i1055(tree_2[983867:982359],tree_2[985376:983868],tree_2[986885:985377],tree_3[656414:654906],tree_3[657923:656415]);
csa_1509 csau_1509_i1056(tree_2[988394:986886],tree_2[989903:988395],tree_2[991412:989904],tree_3[659432:657924],tree_3[660941:659433]);
csa_1509 csau_1509_i1057(tree_2[992921:991413],tree_2[994430:992922],tree_2[995939:994431],tree_3[662450:660942],tree_3[663959:662451]);
csa_1509 csau_1509_i1058(tree_2[997448:995940],tree_2[998957:997449],tree_2[1000466:998958],tree_3[665468:663960],tree_3[666977:665469]);
csa_1509 csau_1509_i1059(tree_2[1001975:1000467],tree_2[1003484:1001976],tree_2[1004993:1003485],tree_3[668486:666978],tree_3[669995:668487]);
csa_1509 csau_1509_i1060(tree_2[1006502:1004994],tree_2[1008011:1006503],tree_2[1009520:1008012],tree_3[671504:669996],tree_3[673013:671505]);
assign tree_3[674522:673014] = tree_2[1011029:1009521];
assign tree_3[676031:674523] = tree_2[1012538:1011030];
// layer-4
csa_1509 csau_1509_i1061(tree_3[1508:0],tree_3[3017:1509],tree_3[4526:3018],tree_4[1508:0],tree_4[3017:1509]);
csa_1509 csau_1509_i1062(tree_3[6035:4527],tree_3[7544:6036],tree_3[9053:7545],tree_4[4526:3018],tree_4[6035:4527]);
csa_1509 csau_1509_i1063(tree_3[10562:9054],tree_3[12071:10563],tree_3[13580:12072],tree_4[7544:6036],tree_4[9053:7545]);
csa_1509 csau_1509_i1064(tree_3[15089:13581],tree_3[16598:15090],tree_3[18107:16599],tree_4[10562:9054],tree_4[12071:10563]);
csa_1509 csau_1509_i1065(tree_3[19616:18108],tree_3[21125:19617],tree_3[22634:21126],tree_4[13580:12072],tree_4[15089:13581]);
csa_1509 csau_1509_i1066(tree_3[24143:22635],tree_3[25652:24144],tree_3[27161:25653],tree_4[16598:15090],tree_4[18107:16599]);
csa_1509 csau_1509_i1067(tree_3[28670:27162],tree_3[30179:28671],tree_3[31688:30180],tree_4[19616:18108],tree_4[21125:19617]);
csa_1509 csau_1509_i1068(tree_3[33197:31689],tree_3[34706:33198],tree_3[36215:34707],tree_4[22634:21126],tree_4[24143:22635]);
csa_1509 csau_1509_i1069(tree_3[37724:36216],tree_3[39233:37725],tree_3[40742:39234],tree_4[25652:24144],tree_4[27161:25653]);
csa_1509 csau_1509_i1070(tree_3[42251:40743],tree_3[43760:42252],tree_3[45269:43761],tree_4[28670:27162],tree_4[30179:28671]);
csa_1509 csau_1509_i1071(tree_3[46778:45270],tree_3[48287:46779],tree_3[49796:48288],tree_4[31688:30180],tree_4[33197:31689]);
csa_1509 csau_1509_i1072(tree_3[51305:49797],tree_3[52814:51306],tree_3[54323:52815],tree_4[34706:33198],tree_4[36215:34707]);
csa_1509 csau_1509_i1073(tree_3[55832:54324],tree_3[57341:55833],tree_3[58850:57342],tree_4[37724:36216],tree_4[39233:37725]);
csa_1509 csau_1509_i1074(tree_3[60359:58851],tree_3[61868:60360],tree_3[63377:61869],tree_4[40742:39234],tree_4[42251:40743]);
csa_1509 csau_1509_i1075(tree_3[64886:63378],tree_3[66395:64887],tree_3[67904:66396],tree_4[43760:42252],tree_4[45269:43761]);
csa_1509 csau_1509_i1076(tree_3[69413:67905],tree_3[70922:69414],tree_3[72431:70923],tree_4[46778:45270],tree_4[48287:46779]);
csa_1509 csau_1509_i1077(tree_3[73940:72432],tree_3[75449:73941],tree_3[76958:75450],tree_4[49796:48288],tree_4[51305:49797]);
csa_1509 csau_1509_i1078(tree_3[78467:76959],tree_3[79976:78468],tree_3[81485:79977],tree_4[52814:51306],tree_4[54323:52815]);
csa_1509 csau_1509_i1079(tree_3[82994:81486],tree_3[84503:82995],tree_3[86012:84504],tree_4[55832:54324],tree_4[57341:55833]);
csa_1509 csau_1509_i1080(tree_3[87521:86013],tree_3[89030:87522],tree_3[90539:89031],tree_4[58850:57342],tree_4[60359:58851]);
csa_1509 csau_1509_i1081(tree_3[92048:90540],tree_3[93557:92049],tree_3[95066:93558],tree_4[61868:60360],tree_4[63377:61869]);
csa_1509 csau_1509_i1082(tree_3[96575:95067],tree_3[98084:96576],tree_3[99593:98085],tree_4[64886:63378],tree_4[66395:64887]);
csa_1509 csau_1509_i1083(tree_3[101102:99594],tree_3[102611:101103],tree_3[104120:102612],tree_4[67904:66396],tree_4[69413:67905]);
csa_1509 csau_1509_i1084(tree_3[105629:104121],tree_3[107138:105630],tree_3[108647:107139],tree_4[70922:69414],tree_4[72431:70923]);
csa_1509 csau_1509_i1085(tree_3[110156:108648],tree_3[111665:110157],tree_3[113174:111666],tree_4[73940:72432],tree_4[75449:73941]);
csa_1509 csau_1509_i1086(tree_3[114683:113175],tree_3[116192:114684],tree_3[117701:116193],tree_4[76958:75450],tree_4[78467:76959]);
csa_1509 csau_1509_i1087(tree_3[119210:117702],tree_3[120719:119211],tree_3[122228:120720],tree_4[79976:78468],tree_4[81485:79977]);
csa_1509 csau_1509_i1088(tree_3[123737:122229],tree_3[125246:123738],tree_3[126755:125247],tree_4[82994:81486],tree_4[84503:82995]);
csa_1509 csau_1509_i1089(tree_3[128264:126756],tree_3[129773:128265],tree_3[131282:129774],tree_4[86012:84504],tree_4[87521:86013]);
csa_1509 csau_1509_i1090(tree_3[132791:131283],tree_3[134300:132792],tree_3[135809:134301],tree_4[89030:87522],tree_4[90539:89031]);
csa_1509 csau_1509_i1091(tree_3[137318:135810],tree_3[138827:137319],tree_3[140336:138828],tree_4[92048:90540],tree_4[93557:92049]);
csa_1509 csau_1509_i1092(tree_3[141845:140337],tree_3[143354:141846],tree_3[144863:143355],tree_4[95066:93558],tree_4[96575:95067]);
csa_1509 csau_1509_i1093(tree_3[146372:144864],tree_3[147881:146373],tree_3[149390:147882],tree_4[98084:96576],tree_4[99593:98085]);
csa_1509 csau_1509_i1094(tree_3[150899:149391],tree_3[152408:150900],tree_3[153917:152409],tree_4[101102:99594],tree_4[102611:101103]);
csa_1509 csau_1509_i1095(tree_3[155426:153918],tree_3[156935:155427],tree_3[158444:156936],tree_4[104120:102612],tree_4[105629:104121]);
csa_1509 csau_1509_i1096(tree_3[159953:158445],tree_3[161462:159954],tree_3[162971:161463],tree_4[107138:105630],tree_4[108647:107139]);
csa_1509 csau_1509_i1097(tree_3[164480:162972],tree_3[165989:164481],tree_3[167498:165990],tree_4[110156:108648],tree_4[111665:110157]);
csa_1509 csau_1509_i1098(tree_3[169007:167499],tree_3[170516:169008],tree_3[172025:170517],tree_4[113174:111666],tree_4[114683:113175]);
csa_1509 csau_1509_i1099(tree_3[173534:172026],tree_3[175043:173535],tree_3[176552:175044],tree_4[116192:114684],tree_4[117701:116193]);
csa_1509 csau_1509_i1100(tree_3[178061:176553],tree_3[179570:178062],tree_3[181079:179571],tree_4[119210:117702],tree_4[120719:119211]);
csa_1509 csau_1509_i1101(tree_3[182588:181080],tree_3[184097:182589],tree_3[185606:184098],tree_4[122228:120720],tree_4[123737:122229]);
csa_1509 csau_1509_i1102(tree_3[187115:185607],tree_3[188624:187116],tree_3[190133:188625],tree_4[125246:123738],tree_4[126755:125247]);
csa_1509 csau_1509_i1103(tree_3[191642:190134],tree_3[193151:191643],tree_3[194660:193152],tree_4[128264:126756],tree_4[129773:128265]);
csa_1509 csau_1509_i1104(tree_3[196169:194661],tree_3[197678:196170],tree_3[199187:197679],tree_4[131282:129774],tree_4[132791:131283]);
csa_1509 csau_1509_i1105(tree_3[200696:199188],tree_3[202205:200697],tree_3[203714:202206],tree_4[134300:132792],tree_4[135809:134301]);
csa_1509 csau_1509_i1106(tree_3[205223:203715],tree_3[206732:205224],tree_3[208241:206733],tree_4[137318:135810],tree_4[138827:137319]);
csa_1509 csau_1509_i1107(tree_3[209750:208242],tree_3[211259:209751],tree_3[212768:211260],tree_4[140336:138828],tree_4[141845:140337]);
csa_1509 csau_1509_i1108(tree_3[214277:212769],tree_3[215786:214278],tree_3[217295:215787],tree_4[143354:141846],tree_4[144863:143355]);
csa_1509 csau_1509_i1109(tree_3[218804:217296],tree_3[220313:218805],tree_3[221822:220314],tree_4[146372:144864],tree_4[147881:146373]);
csa_1509 csau_1509_i1110(tree_3[223331:221823],tree_3[224840:223332],tree_3[226349:224841],tree_4[149390:147882],tree_4[150899:149391]);
csa_1509 csau_1509_i1111(tree_3[227858:226350],tree_3[229367:227859],tree_3[230876:229368],tree_4[152408:150900],tree_4[153917:152409]);
csa_1509 csau_1509_i1112(tree_3[232385:230877],tree_3[233894:232386],tree_3[235403:233895],tree_4[155426:153918],tree_4[156935:155427]);
csa_1509 csau_1509_i1113(tree_3[236912:235404],tree_3[238421:236913],tree_3[239930:238422],tree_4[158444:156936],tree_4[159953:158445]);
csa_1509 csau_1509_i1114(tree_3[241439:239931],tree_3[242948:241440],tree_3[244457:242949],tree_4[161462:159954],tree_4[162971:161463]);
csa_1509 csau_1509_i1115(tree_3[245966:244458],tree_3[247475:245967],tree_3[248984:247476],tree_4[164480:162972],tree_4[165989:164481]);
csa_1509 csau_1509_i1116(tree_3[250493:248985],tree_3[252002:250494],tree_3[253511:252003],tree_4[167498:165990],tree_4[169007:167499]);
csa_1509 csau_1509_i1117(tree_3[255020:253512],tree_3[256529:255021],tree_3[258038:256530],tree_4[170516:169008],tree_4[172025:170517]);
csa_1509 csau_1509_i1118(tree_3[259547:258039],tree_3[261056:259548],tree_3[262565:261057],tree_4[173534:172026],tree_4[175043:173535]);
csa_1509 csau_1509_i1119(tree_3[264074:262566],tree_3[265583:264075],tree_3[267092:265584],tree_4[176552:175044],tree_4[178061:176553]);
csa_1509 csau_1509_i1120(tree_3[268601:267093],tree_3[270110:268602],tree_3[271619:270111],tree_4[179570:178062],tree_4[181079:179571]);
csa_1509 csau_1509_i1121(tree_3[273128:271620],tree_3[274637:273129],tree_3[276146:274638],tree_4[182588:181080],tree_4[184097:182589]);
csa_1509 csau_1509_i1122(tree_3[277655:276147],tree_3[279164:277656],tree_3[280673:279165],tree_4[185606:184098],tree_4[187115:185607]);
csa_1509 csau_1509_i1123(tree_3[282182:280674],tree_3[283691:282183],tree_3[285200:283692],tree_4[188624:187116],tree_4[190133:188625]);
csa_1509 csau_1509_i1124(tree_3[286709:285201],tree_3[288218:286710],tree_3[289727:288219],tree_4[191642:190134],tree_4[193151:191643]);
csa_1509 csau_1509_i1125(tree_3[291236:289728],tree_3[292745:291237],tree_3[294254:292746],tree_4[194660:193152],tree_4[196169:194661]);
csa_1509 csau_1509_i1126(tree_3[295763:294255],tree_3[297272:295764],tree_3[298781:297273],tree_4[197678:196170],tree_4[199187:197679]);
csa_1509 csau_1509_i1127(tree_3[300290:298782],tree_3[301799:300291],tree_3[303308:301800],tree_4[200696:199188],tree_4[202205:200697]);
csa_1509 csau_1509_i1128(tree_3[304817:303309],tree_3[306326:304818],tree_3[307835:306327],tree_4[203714:202206],tree_4[205223:203715]);
csa_1509 csau_1509_i1129(tree_3[309344:307836],tree_3[310853:309345],tree_3[312362:310854],tree_4[206732:205224],tree_4[208241:206733]);
csa_1509 csau_1509_i1130(tree_3[313871:312363],tree_3[315380:313872],tree_3[316889:315381],tree_4[209750:208242],tree_4[211259:209751]);
csa_1509 csau_1509_i1131(tree_3[318398:316890],tree_3[319907:318399],tree_3[321416:319908],tree_4[212768:211260],tree_4[214277:212769]);
csa_1509 csau_1509_i1132(tree_3[322925:321417],tree_3[324434:322926],tree_3[325943:324435],tree_4[215786:214278],tree_4[217295:215787]);
csa_1509 csau_1509_i1133(tree_3[327452:325944],tree_3[328961:327453],tree_3[330470:328962],tree_4[218804:217296],tree_4[220313:218805]);
csa_1509 csau_1509_i1134(tree_3[331979:330471],tree_3[333488:331980],tree_3[334997:333489],tree_4[221822:220314],tree_4[223331:221823]);
csa_1509 csau_1509_i1135(tree_3[336506:334998],tree_3[338015:336507],tree_3[339524:338016],tree_4[224840:223332],tree_4[226349:224841]);
csa_1509 csau_1509_i1136(tree_3[341033:339525],tree_3[342542:341034],tree_3[344051:342543],tree_4[227858:226350],tree_4[229367:227859]);
csa_1509 csau_1509_i1137(tree_3[345560:344052],tree_3[347069:345561],tree_3[348578:347070],tree_4[230876:229368],tree_4[232385:230877]);
csa_1509 csau_1509_i1138(tree_3[350087:348579],tree_3[351596:350088],tree_3[353105:351597],tree_4[233894:232386],tree_4[235403:233895]);
csa_1509 csau_1509_i1139(tree_3[354614:353106],tree_3[356123:354615],tree_3[357632:356124],tree_4[236912:235404],tree_4[238421:236913]);
csa_1509 csau_1509_i1140(tree_3[359141:357633],tree_3[360650:359142],tree_3[362159:360651],tree_4[239930:238422],tree_4[241439:239931]);
csa_1509 csau_1509_i1141(tree_3[363668:362160],tree_3[365177:363669],tree_3[366686:365178],tree_4[242948:241440],tree_4[244457:242949]);
csa_1509 csau_1509_i1142(tree_3[368195:366687],tree_3[369704:368196],tree_3[371213:369705],tree_4[245966:244458],tree_4[247475:245967]);
csa_1509 csau_1509_i1143(tree_3[372722:371214],tree_3[374231:372723],tree_3[375740:374232],tree_4[248984:247476],tree_4[250493:248985]);
csa_1509 csau_1509_i1144(tree_3[377249:375741],tree_3[378758:377250],tree_3[380267:378759],tree_4[252002:250494],tree_4[253511:252003]);
csa_1509 csau_1509_i1145(tree_3[381776:380268],tree_3[383285:381777],tree_3[384794:383286],tree_4[255020:253512],tree_4[256529:255021]);
csa_1509 csau_1509_i1146(tree_3[386303:384795],tree_3[387812:386304],tree_3[389321:387813],tree_4[258038:256530],tree_4[259547:258039]);
csa_1509 csau_1509_i1147(tree_3[390830:389322],tree_3[392339:390831],tree_3[393848:392340],tree_4[261056:259548],tree_4[262565:261057]);
csa_1509 csau_1509_i1148(tree_3[395357:393849],tree_3[396866:395358],tree_3[398375:396867],tree_4[264074:262566],tree_4[265583:264075]);
csa_1509 csau_1509_i1149(tree_3[399884:398376],tree_3[401393:399885],tree_3[402902:401394],tree_4[267092:265584],tree_4[268601:267093]);
csa_1509 csau_1509_i1150(tree_3[404411:402903],tree_3[405920:404412],tree_3[407429:405921],tree_4[270110:268602],tree_4[271619:270111]);
csa_1509 csau_1509_i1151(tree_3[408938:407430],tree_3[410447:408939],tree_3[411956:410448],tree_4[273128:271620],tree_4[274637:273129]);
csa_1509 csau_1509_i1152(tree_3[413465:411957],tree_3[414974:413466],tree_3[416483:414975],tree_4[276146:274638],tree_4[277655:276147]);
csa_1509 csau_1509_i1153(tree_3[417992:416484],tree_3[419501:417993],tree_3[421010:419502],tree_4[279164:277656],tree_4[280673:279165]);
csa_1509 csau_1509_i1154(tree_3[422519:421011],tree_3[424028:422520],tree_3[425537:424029],tree_4[282182:280674],tree_4[283691:282183]);
csa_1509 csau_1509_i1155(tree_3[427046:425538],tree_3[428555:427047],tree_3[430064:428556],tree_4[285200:283692],tree_4[286709:285201]);
csa_1509 csau_1509_i1156(tree_3[431573:430065],tree_3[433082:431574],tree_3[434591:433083],tree_4[288218:286710],tree_4[289727:288219]);
csa_1509 csau_1509_i1157(tree_3[436100:434592],tree_3[437609:436101],tree_3[439118:437610],tree_4[291236:289728],tree_4[292745:291237]);
csa_1509 csau_1509_i1158(tree_3[440627:439119],tree_3[442136:440628],tree_3[443645:442137],tree_4[294254:292746],tree_4[295763:294255]);
csa_1509 csau_1509_i1159(tree_3[445154:443646],tree_3[446663:445155],tree_3[448172:446664],tree_4[297272:295764],tree_4[298781:297273]);
csa_1509 csau_1509_i1160(tree_3[449681:448173],tree_3[451190:449682],tree_3[452699:451191],tree_4[300290:298782],tree_4[301799:300291]);
csa_1509 csau_1509_i1161(tree_3[454208:452700],tree_3[455717:454209],tree_3[457226:455718],tree_4[303308:301800],tree_4[304817:303309]);
csa_1509 csau_1509_i1162(tree_3[458735:457227],tree_3[460244:458736],tree_3[461753:460245],tree_4[306326:304818],tree_4[307835:306327]);
csa_1509 csau_1509_i1163(tree_3[463262:461754],tree_3[464771:463263],tree_3[466280:464772],tree_4[309344:307836],tree_4[310853:309345]);
csa_1509 csau_1509_i1164(tree_3[467789:466281],tree_3[469298:467790],tree_3[470807:469299],tree_4[312362:310854],tree_4[313871:312363]);
csa_1509 csau_1509_i1165(tree_3[472316:470808],tree_3[473825:472317],tree_3[475334:473826],tree_4[315380:313872],tree_4[316889:315381]);
csa_1509 csau_1509_i1166(tree_3[476843:475335],tree_3[478352:476844],tree_3[479861:478353],tree_4[318398:316890],tree_4[319907:318399]);
csa_1509 csau_1509_i1167(tree_3[481370:479862],tree_3[482879:481371],tree_3[484388:482880],tree_4[321416:319908],tree_4[322925:321417]);
csa_1509 csau_1509_i1168(tree_3[485897:484389],tree_3[487406:485898],tree_3[488915:487407],tree_4[324434:322926],tree_4[325943:324435]);
csa_1509 csau_1509_i1169(tree_3[490424:488916],tree_3[491933:490425],tree_3[493442:491934],tree_4[327452:325944],tree_4[328961:327453]);
csa_1509 csau_1509_i1170(tree_3[494951:493443],tree_3[496460:494952],tree_3[497969:496461],tree_4[330470:328962],tree_4[331979:330471]);
csa_1509 csau_1509_i1171(tree_3[499478:497970],tree_3[500987:499479],tree_3[502496:500988],tree_4[333488:331980],tree_4[334997:333489]);
csa_1509 csau_1509_i1172(tree_3[504005:502497],tree_3[505514:504006],tree_3[507023:505515],tree_4[336506:334998],tree_4[338015:336507]);
csa_1509 csau_1509_i1173(tree_3[508532:507024],tree_3[510041:508533],tree_3[511550:510042],tree_4[339524:338016],tree_4[341033:339525]);
csa_1509 csau_1509_i1174(tree_3[513059:511551],tree_3[514568:513060],tree_3[516077:514569],tree_4[342542:341034],tree_4[344051:342543]);
csa_1509 csau_1509_i1175(tree_3[517586:516078],tree_3[519095:517587],tree_3[520604:519096],tree_4[345560:344052],tree_4[347069:345561]);
csa_1509 csau_1509_i1176(tree_3[522113:520605],tree_3[523622:522114],tree_3[525131:523623],tree_4[348578:347070],tree_4[350087:348579]);
csa_1509 csau_1509_i1177(tree_3[526640:525132],tree_3[528149:526641],tree_3[529658:528150],tree_4[351596:350088],tree_4[353105:351597]);
csa_1509 csau_1509_i1178(tree_3[531167:529659],tree_3[532676:531168],tree_3[534185:532677],tree_4[354614:353106],tree_4[356123:354615]);
csa_1509 csau_1509_i1179(tree_3[535694:534186],tree_3[537203:535695],tree_3[538712:537204],tree_4[357632:356124],tree_4[359141:357633]);
csa_1509 csau_1509_i1180(tree_3[540221:538713],tree_3[541730:540222],tree_3[543239:541731],tree_4[360650:359142],tree_4[362159:360651]);
csa_1509 csau_1509_i1181(tree_3[544748:543240],tree_3[546257:544749],tree_3[547766:546258],tree_4[363668:362160],tree_4[365177:363669]);
csa_1509 csau_1509_i1182(tree_3[549275:547767],tree_3[550784:549276],tree_3[552293:550785],tree_4[366686:365178],tree_4[368195:366687]);
csa_1509 csau_1509_i1183(tree_3[553802:552294],tree_3[555311:553803],tree_3[556820:555312],tree_4[369704:368196],tree_4[371213:369705]);
csa_1509 csau_1509_i1184(tree_3[558329:556821],tree_3[559838:558330],tree_3[561347:559839],tree_4[372722:371214],tree_4[374231:372723]);
csa_1509 csau_1509_i1185(tree_3[562856:561348],tree_3[564365:562857],tree_3[565874:564366],tree_4[375740:374232],tree_4[377249:375741]);
csa_1509 csau_1509_i1186(tree_3[567383:565875],tree_3[568892:567384],tree_3[570401:568893],tree_4[378758:377250],tree_4[380267:378759]);
csa_1509 csau_1509_i1187(tree_3[571910:570402],tree_3[573419:571911],tree_3[574928:573420],tree_4[381776:380268],tree_4[383285:381777]);
csa_1509 csau_1509_i1188(tree_3[576437:574929],tree_3[577946:576438],tree_3[579455:577947],tree_4[384794:383286],tree_4[386303:384795]);
csa_1509 csau_1509_i1189(tree_3[580964:579456],tree_3[582473:580965],tree_3[583982:582474],tree_4[387812:386304],tree_4[389321:387813]);
csa_1509 csau_1509_i1190(tree_3[585491:583983],tree_3[587000:585492],tree_3[588509:587001],tree_4[390830:389322],tree_4[392339:390831]);
csa_1509 csau_1509_i1191(tree_3[590018:588510],tree_3[591527:590019],tree_3[593036:591528],tree_4[393848:392340],tree_4[395357:393849]);
csa_1509 csau_1509_i1192(tree_3[594545:593037],tree_3[596054:594546],tree_3[597563:596055],tree_4[396866:395358],tree_4[398375:396867]);
csa_1509 csau_1509_i1193(tree_3[599072:597564],tree_3[600581:599073],tree_3[602090:600582],tree_4[399884:398376],tree_4[401393:399885]);
csa_1509 csau_1509_i1194(tree_3[603599:602091],tree_3[605108:603600],tree_3[606617:605109],tree_4[402902:401394],tree_4[404411:402903]);
csa_1509 csau_1509_i1195(tree_3[608126:606618],tree_3[609635:608127],tree_3[611144:609636],tree_4[405920:404412],tree_4[407429:405921]);
csa_1509 csau_1509_i1196(tree_3[612653:611145],tree_3[614162:612654],tree_3[615671:614163],tree_4[408938:407430],tree_4[410447:408939]);
csa_1509 csau_1509_i1197(tree_3[617180:615672],tree_3[618689:617181],tree_3[620198:618690],tree_4[411956:410448],tree_4[413465:411957]);
csa_1509 csau_1509_i1198(tree_3[621707:620199],tree_3[623216:621708],tree_3[624725:623217],tree_4[414974:413466],tree_4[416483:414975]);
csa_1509 csau_1509_i1199(tree_3[626234:624726],tree_3[627743:626235],tree_3[629252:627744],tree_4[417992:416484],tree_4[419501:417993]);
csa_1509 csau_1509_i1200(tree_3[630761:629253],tree_3[632270:630762],tree_3[633779:632271],tree_4[421010:419502],tree_4[422519:421011]);
csa_1509 csau_1509_i1201(tree_3[635288:633780],tree_3[636797:635289],tree_3[638306:636798],tree_4[424028:422520],tree_4[425537:424029]);
csa_1509 csau_1509_i1202(tree_3[639815:638307],tree_3[641324:639816],tree_3[642833:641325],tree_4[427046:425538],tree_4[428555:427047]);
csa_1509 csau_1509_i1203(tree_3[644342:642834],tree_3[645851:644343],tree_3[647360:645852],tree_4[430064:428556],tree_4[431573:430065]);
csa_1509 csau_1509_i1204(tree_3[648869:647361],tree_3[650378:648870],tree_3[651887:650379],tree_4[433082:431574],tree_4[434591:433083]);
csa_1509 csau_1509_i1205(tree_3[653396:651888],tree_3[654905:653397],tree_3[656414:654906],tree_4[436100:434592],tree_4[437609:436101]);
csa_1509 csau_1509_i1206(tree_3[657923:656415],tree_3[659432:657924],tree_3[660941:659433],tree_4[439118:437610],tree_4[440627:439119]);
csa_1509 csau_1509_i1207(tree_3[662450:660942],tree_3[663959:662451],tree_3[665468:663960],tree_4[442136:440628],tree_4[443645:442137]);
csa_1509 csau_1509_i1208(tree_3[666977:665469],tree_3[668486:666978],tree_3[669995:668487],tree_4[445154:443646],tree_4[446663:445155]);
csa_1509 csau_1509_i1209(tree_3[671504:669996],tree_3[673013:671505],tree_3[674522:673014],tree_4[448172:446664],tree_4[449681:448173]);
assign tree_4[451190:449682] = tree_3[676031:674523];
// layer-5
csa_1509 csau_1509_i1210(tree_4[1508:0],tree_4[3017:1509],tree_4[4526:3018],tree_5[1508:0],tree_5[3017:1509]);
csa_1509 csau_1509_i1211(tree_4[6035:4527],tree_4[7544:6036],tree_4[9053:7545],tree_5[4526:3018],tree_5[6035:4527]);
csa_1509 csau_1509_i1212(tree_4[10562:9054],tree_4[12071:10563],tree_4[13580:12072],tree_5[7544:6036],tree_5[9053:7545]);
csa_1509 csau_1509_i1213(tree_4[15089:13581],tree_4[16598:15090],tree_4[18107:16599],tree_5[10562:9054],tree_5[12071:10563]);
csa_1509 csau_1509_i1214(tree_4[19616:18108],tree_4[21125:19617],tree_4[22634:21126],tree_5[13580:12072],tree_5[15089:13581]);
csa_1509 csau_1509_i1215(tree_4[24143:22635],tree_4[25652:24144],tree_4[27161:25653],tree_5[16598:15090],tree_5[18107:16599]);
csa_1509 csau_1509_i1216(tree_4[28670:27162],tree_4[30179:28671],tree_4[31688:30180],tree_5[19616:18108],tree_5[21125:19617]);
csa_1509 csau_1509_i1217(tree_4[33197:31689],tree_4[34706:33198],tree_4[36215:34707],tree_5[22634:21126],tree_5[24143:22635]);
csa_1509 csau_1509_i1218(tree_4[37724:36216],tree_4[39233:37725],tree_4[40742:39234],tree_5[25652:24144],tree_5[27161:25653]);
csa_1509 csau_1509_i1219(tree_4[42251:40743],tree_4[43760:42252],tree_4[45269:43761],tree_5[28670:27162],tree_5[30179:28671]);
csa_1509 csau_1509_i1220(tree_4[46778:45270],tree_4[48287:46779],tree_4[49796:48288],tree_5[31688:30180],tree_5[33197:31689]);
csa_1509 csau_1509_i1221(tree_4[51305:49797],tree_4[52814:51306],tree_4[54323:52815],tree_5[34706:33198],tree_5[36215:34707]);
csa_1509 csau_1509_i1222(tree_4[55832:54324],tree_4[57341:55833],tree_4[58850:57342],tree_5[37724:36216],tree_5[39233:37725]);
csa_1509 csau_1509_i1223(tree_4[60359:58851],tree_4[61868:60360],tree_4[63377:61869],tree_5[40742:39234],tree_5[42251:40743]);
csa_1509 csau_1509_i1224(tree_4[64886:63378],tree_4[66395:64887],tree_4[67904:66396],tree_5[43760:42252],tree_5[45269:43761]);
csa_1509 csau_1509_i1225(tree_4[69413:67905],tree_4[70922:69414],tree_4[72431:70923],tree_5[46778:45270],tree_5[48287:46779]);
csa_1509 csau_1509_i1226(tree_4[73940:72432],tree_4[75449:73941],tree_4[76958:75450],tree_5[49796:48288],tree_5[51305:49797]);
csa_1509 csau_1509_i1227(tree_4[78467:76959],tree_4[79976:78468],tree_4[81485:79977],tree_5[52814:51306],tree_5[54323:52815]);
csa_1509 csau_1509_i1228(tree_4[82994:81486],tree_4[84503:82995],tree_4[86012:84504],tree_5[55832:54324],tree_5[57341:55833]);
csa_1509 csau_1509_i1229(tree_4[87521:86013],tree_4[89030:87522],tree_4[90539:89031],tree_5[58850:57342],tree_5[60359:58851]);
csa_1509 csau_1509_i1230(tree_4[92048:90540],tree_4[93557:92049],tree_4[95066:93558],tree_5[61868:60360],tree_5[63377:61869]);
csa_1509 csau_1509_i1231(tree_4[96575:95067],tree_4[98084:96576],tree_4[99593:98085],tree_5[64886:63378],tree_5[66395:64887]);
csa_1509 csau_1509_i1232(tree_4[101102:99594],tree_4[102611:101103],tree_4[104120:102612],tree_5[67904:66396],tree_5[69413:67905]);
csa_1509 csau_1509_i1233(tree_4[105629:104121],tree_4[107138:105630],tree_4[108647:107139],tree_5[70922:69414],tree_5[72431:70923]);
csa_1509 csau_1509_i1234(tree_4[110156:108648],tree_4[111665:110157],tree_4[113174:111666],tree_5[73940:72432],tree_5[75449:73941]);
csa_1509 csau_1509_i1235(tree_4[114683:113175],tree_4[116192:114684],tree_4[117701:116193],tree_5[76958:75450],tree_5[78467:76959]);
csa_1509 csau_1509_i1236(tree_4[119210:117702],tree_4[120719:119211],tree_4[122228:120720],tree_5[79976:78468],tree_5[81485:79977]);
csa_1509 csau_1509_i1237(tree_4[123737:122229],tree_4[125246:123738],tree_4[126755:125247],tree_5[82994:81486],tree_5[84503:82995]);
csa_1509 csau_1509_i1238(tree_4[128264:126756],tree_4[129773:128265],tree_4[131282:129774],tree_5[86012:84504],tree_5[87521:86013]);
csa_1509 csau_1509_i1239(tree_4[132791:131283],tree_4[134300:132792],tree_4[135809:134301],tree_5[89030:87522],tree_5[90539:89031]);
csa_1509 csau_1509_i1240(tree_4[137318:135810],tree_4[138827:137319],tree_4[140336:138828],tree_5[92048:90540],tree_5[93557:92049]);
csa_1509 csau_1509_i1241(tree_4[141845:140337],tree_4[143354:141846],tree_4[144863:143355],tree_5[95066:93558],tree_5[96575:95067]);
csa_1509 csau_1509_i1242(tree_4[146372:144864],tree_4[147881:146373],tree_4[149390:147882],tree_5[98084:96576],tree_5[99593:98085]);
csa_1509 csau_1509_i1243(tree_4[150899:149391],tree_4[152408:150900],tree_4[153917:152409],tree_5[101102:99594],tree_5[102611:101103]);
csa_1509 csau_1509_i1244(tree_4[155426:153918],tree_4[156935:155427],tree_4[158444:156936],tree_5[104120:102612],tree_5[105629:104121]);
csa_1509 csau_1509_i1245(tree_4[159953:158445],tree_4[161462:159954],tree_4[162971:161463],tree_5[107138:105630],tree_5[108647:107139]);
csa_1509 csau_1509_i1246(tree_4[164480:162972],tree_4[165989:164481],tree_4[167498:165990],tree_5[110156:108648],tree_5[111665:110157]);
csa_1509 csau_1509_i1247(tree_4[169007:167499],tree_4[170516:169008],tree_4[172025:170517],tree_5[113174:111666],tree_5[114683:113175]);
csa_1509 csau_1509_i1248(tree_4[173534:172026],tree_4[175043:173535],tree_4[176552:175044],tree_5[116192:114684],tree_5[117701:116193]);
csa_1509 csau_1509_i1249(tree_4[178061:176553],tree_4[179570:178062],tree_4[181079:179571],tree_5[119210:117702],tree_5[120719:119211]);
csa_1509 csau_1509_i1250(tree_4[182588:181080],tree_4[184097:182589],tree_4[185606:184098],tree_5[122228:120720],tree_5[123737:122229]);
csa_1509 csau_1509_i1251(tree_4[187115:185607],tree_4[188624:187116],tree_4[190133:188625],tree_5[125246:123738],tree_5[126755:125247]);
csa_1509 csau_1509_i1252(tree_4[191642:190134],tree_4[193151:191643],tree_4[194660:193152],tree_5[128264:126756],tree_5[129773:128265]);
csa_1509 csau_1509_i1253(tree_4[196169:194661],tree_4[197678:196170],tree_4[199187:197679],tree_5[131282:129774],tree_5[132791:131283]);
csa_1509 csau_1509_i1254(tree_4[200696:199188],tree_4[202205:200697],tree_4[203714:202206],tree_5[134300:132792],tree_5[135809:134301]);
csa_1509 csau_1509_i1255(tree_4[205223:203715],tree_4[206732:205224],tree_4[208241:206733],tree_5[137318:135810],tree_5[138827:137319]);
csa_1509 csau_1509_i1256(tree_4[209750:208242],tree_4[211259:209751],tree_4[212768:211260],tree_5[140336:138828],tree_5[141845:140337]);
csa_1509 csau_1509_i1257(tree_4[214277:212769],tree_4[215786:214278],tree_4[217295:215787],tree_5[143354:141846],tree_5[144863:143355]);
csa_1509 csau_1509_i1258(tree_4[218804:217296],tree_4[220313:218805],tree_4[221822:220314],tree_5[146372:144864],tree_5[147881:146373]);
csa_1509 csau_1509_i1259(tree_4[223331:221823],tree_4[224840:223332],tree_4[226349:224841],tree_5[149390:147882],tree_5[150899:149391]);
csa_1509 csau_1509_i1260(tree_4[227858:226350],tree_4[229367:227859],tree_4[230876:229368],tree_5[152408:150900],tree_5[153917:152409]);
csa_1509 csau_1509_i1261(tree_4[232385:230877],tree_4[233894:232386],tree_4[235403:233895],tree_5[155426:153918],tree_5[156935:155427]);
csa_1509 csau_1509_i1262(tree_4[236912:235404],tree_4[238421:236913],tree_4[239930:238422],tree_5[158444:156936],tree_5[159953:158445]);
csa_1509 csau_1509_i1263(tree_4[241439:239931],tree_4[242948:241440],tree_4[244457:242949],tree_5[161462:159954],tree_5[162971:161463]);
csa_1509 csau_1509_i1264(tree_4[245966:244458],tree_4[247475:245967],tree_4[248984:247476],tree_5[164480:162972],tree_5[165989:164481]);
csa_1509 csau_1509_i1265(tree_4[250493:248985],tree_4[252002:250494],tree_4[253511:252003],tree_5[167498:165990],tree_5[169007:167499]);
csa_1509 csau_1509_i1266(tree_4[255020:253512],tree_4[256529:255021],tree_4[258038:256530],tree_5[170516:169008],tree_5[172025:170517]);
csa_1509 csau_1509_i1267(tree_4[259547:258039],tree_4[261056:259548],tree_4[262565:261057],tree_5[173534:172026],tree_5[175043:173535]);
csa_1509 csau_1509_i1268(tree_4[264074:262566],tree_4[265583:264075],tree_4[267092:265584],tree_5[176552:175044],tree_5[178061:176553]);
csa_1509 csau_1509_i1269(tree_4[268601:267093],tree_4[270110:268602],tree_4[271619:270111],tree_5[179570:178062],tree_5[181079:179571]);
csa_1509 csau_1509_i1270(tree_4[273128:271620],tree_4[274637:273129],tree_4[276146:274638],tree_5[182588:181080],tree_5[184097:182589]);
csa_1509 csau_1509_i1271(tree_4[277655:276147],tree_4[279164:277656],tree_4[280673:279165],tree_5[185606:184098],tree_5[187115:185607]);
csa_1509 csau_1509_i1272(tree_4[282182:280674],tree_4[283691:282183],tree_4[285200:283692],tree_5[188624:187116],tree_5[190133:188625]);
csa_1509 csau_1509_i1273(tree_4[286709:285201],tree_4[288218:286710],tree_4[289727:288219],tree_5[191642:190134],tree_5[193151:191643]);
csa_1509 csau_1509_i1274(tree_4[291236:289728],tree_4[292745:291237],tree_4[294254:292746],tree_5[194660:193152],tree_5[196169:194661]);
csa_1509 csau_1509_i1275(tree_4[295763:294255],tree_4[297272:295764],tree_4[298781:297273],tree_5[197678:196170],tree_5[199187:197679]);
csa_1509 csau_1509_i1276(tree_4[300290:298782],tree_4[301799:300291],tree_4[303308:301800],tree_5[200696:199188],tree_5[202205:200697]);
csa_1509 csau_1509_i1277(tree_4[304817:303309],tree_4[306326:304818],tree_4[307835:306327],tree_5[203714:202206],tree_5[205223:203715]);
csa_1509 csau_1509_i1278(tree_4[309344:307836],tree_4[310853:309345],tree_4[312362:310854],tree_5[206732:205224],tree_5[208241:206733]);
csa_1509 csau_1509_i1279(tree_4[313871:312363],tree_4[315380:313872],tree_4[316889:315381],tree_5[209750:208242],tree_5[211259:209751]);
csa_1509 csau_1509_i1280(tree_4[318398:316890],tree_4[319907:318399],tree_4[321416:319908],tree_5[212768:211260],tree_5[214277:212769]);
csa_1509 csau_1509_i1281(tree_4[322925:321417],tree_4[324434:322926],tree_4[325943:324435],tree_5[215786:214278],tree_5[217295:215787]);
csa_1509 csau_1509_i1282(tree_4[327452:325944],tree_4[328961:327453],tree_4[330470:328962],tree_5[218804:217296],tree_5[220313:218805]);
csa_1509 csau_1509_i1283(tree_4[331979:330471],tree_4[333488:331980],tree_4[334997:333489],tree_5[221822:220314],tree_5[223331:221823]);
csa_1509 csau_1509_i1284(tree_4[336506:334998],tree_4[338015:336507],tree_4[339524:338016],tree_5[224840:223332],tree_5[226349:224841]);
csa_1509 csau_1509_i1285(tree_4[341033:339525],tree_4[342542:341034],tree_4[344051:342543],tree_5[227858:226350],tree_5[229367:227859]);
csa_1509 csau_1509_i1286(tree_4[345560:344052],tree_4[347069:345561],tree_4[348578:347070],tree_5[230876:229368],tree_5[232385:230877]);
csa_1509 csau_1509_i1287(tree_4[350087:348579],tree_4[351596:350088],tree_4[353105:351597],tree_5[233894:232386],tree_5[235403:233895]);
csa_1509 csau_1509_i1288(tree_4[354614:353106],tree_4[356123:354615],tree_4[357632:356124],tree_5[236912:235404],tree_5[238421:236913]);
csa_1509 csau_1509_i1289(tree_4[359141:357633],tree_4[360650:359142],tree_4[362159:360651],tree_5[239930:238422],tree_5[241439:239931]);
csa_1509 csau_1509_i1290(tree_4[363668:362160],tree_4[365177:363669],tree_4[366686:365178],tree_5[242948:241440],tree_5[244457:242949]);
csa_1509 csau_1509_i1291(tree_4[368195:366687],tree_4[369704:368196],tree_4[371213:369705],tree_5[245966:244458],tree_5[247475:245967]);
csa_1509 csau_1509_i1292(tree_4[372722:371214],tree_4[374231:372723],tree_4[375740:374232],tree_5[248984:247476],tree_5[250493:248985]);
csa_1509 csau_1509_i1293(tree_4[377249:375741],tree_4[378758:377250],tree_4[380267:378759],tree_5[252002:250494],tree_5[253511:252003]);
csa_1509 csau_1509_i1294(tree_4[381776:380268],tree_4[383285:381777],tree_4[384794:383286],tree_5[255020:253512],tree_5[256529:255021]);
csa_1509 csau_1509_i1295(tree_4[386303:384795],tree_4[387812:386304],tree_4[389321:387813],tree_5[258038:256530],tree_5[259547:258039]);
csa_1509 csau_1509_i1296(tree_4[390830:389322],tree_4[392339:390831],tree_4[393848:392340],tree_5[261056:259548],tree_5[262565:261057]);
csa_1509 csau_1509_i1297(tree_4[395357:393849],tree_4[396866:395358],tree_4[398375:396867],tree_5[264074:262566],tree_5[265583:264075]);
csa_1509 csau_1509_i1298(tree_4[399884:398376],tree_4[401393:399885],tree_4[402902:401394],tree_5[267092:265584],tree_5[268601:267093]);
csa_1509 csau_1509_i1299(tree_4[404411:402903],tree_4[405920:404412],tree_4[407429:405921],tree_5[270110:268602],tree_5[271619:270111]);
csa_1509 csau_1509_i1300(tree_4[408938:407430],tree_4[410447:408939],tree_4[411956:410448],tree_5[273128:271620],tree_5[274637:273129]);
csa_1509 csau_1509_i1301(tree_4[413465:411957],tree_4[414974:413466],tree_4[416483:414975],tree_5[276146:274638],tree_5[277655:276147]);
csa_1509 csau_1509_i1302(tree_4[417992:416484],tree_4[419501:417993],tree_4[421010:419502],tree_5[279164:277656],tree_5[280673:279165]);
csa_1509 csau_1509_i1303(tree_4[422519:421011],tree_4[424028:422520],tree_4[425537:424029],tree_5[282182:280674],tree_5[283691:282183]);
csa_1509 csau_1509_i1304(tree_4[427046:425538],tree_4[428555:427047],tree_4[430064:428556],tree_5[285200:283692],tree_5[286709:285201]);
csa_1509 csau_1509_i1305(tree_4[431573:430065],tree_4[433082:431574],tree_4[434591:433083],tree_5[288218:286710],tree_5[289727:288219]);
csa_1509 csau_1509_i1306(tree_4[436100:434592],tree_4[437609:436101],tree_4[439118:437610],tree_5[291236:289728],tree_5[292745:291237]);
csa_1509 csau_1509_i1307(tree_4[440627:439119],tree_4[442136:440628],tree_4[443645:442137],tree_5[294254:292746],tree_5[295763:294255]);
csa_1509 csau_1509_i1308(tree_4[445154:443646],tree_4[446663:445155],tree_4[448172:446664],tree_5[297272:295764],tree_5[298781:297273]);
assign tree_5[300290:298782] = tree_4[449681:448173];
assign tree_5[301799:300291] = tree_4[451190:449682];
// layer-6
csa_1509 csau_1509_i1309(tree_5[1508:0],tree_5[3017:1509],tree_5[4526:3018],tree_6[1508:0],tree_6[3017:1509]);
csa_1509 csau_1509_i1310(tree_5[6035:4527],tree_5[7544:6036],tree_5[9053:7545],tree_6[4526:3018],tree_6[6035:4527]);
csa_1509 csau_1509_i1311(tree_5[10562:9054],tree_5[12071:10563],tree_5[13580:12072],tree_6[7544:6036],tree_6[9053:7545]);
csa_1509 csau_1509_i1312(tree_5[15089:13581],tree_5[16598:15090],tree_5[18107:16599],tree_6[10562:9054],tree_6[12071:10563]);
csa_1509 csau_1509_i1313(tree_5[19616:18108],tree_5[21125:19617],tree_5[22634:21126],tree_6[13580:12072],tree_6[15089:13581]);
csa_1509 csau_1509_i1314(tree_5[24143:22635],tree_5[25652:24144],tree_5[27161:25653],tree_6[16598:15090],tree_6[18107:16599]);
csa_1509 csau_1509_i1315(tree_5[28670:27162],tree_5[30179:28671],tree_5[31688:30180],tree_6[19616:18108],tree_6[21125:19617]);
csa_1509 csau_1509_i1316(tree_5[33197:31689],tree_5[34706:33198],tree_5[36215:34707],tree_6[22634:21126],tree_6[24143:22635]);
csa_1509 csau_1509_i1317(tree_5[37724:36216],tree_5[39233:37725],tree_5[40742:39234],tree_6[25652:24144],tree_6[27161:25653]);
csa_1509 csau_1509_i1318(tree_5[42251:40743],tree_5[43760:42252],tree_5[45269:43761],tree_6[28670:27162],tree_6[30179:28671]);
csa_1509 csau_1509_i1319(tree_5[46778:45270],tree_5[48287:46779],tree_5[49796:48288],tree_6[31688:30180],tree_6[33197:31689]);
csa_1509 csau_1509_i1320(tree_5[51305:49797],tree_5[52814:51306],tree_5[54323:52815],tree_6[34706:33198],tree_6[36215:34707]);
csa_1509 csau_1509_i1321(tree_5[55832:54324],tree_5[57341:55833],tree_5[58850:57342],tree_6[37724:36216],tree_6[39233:37725]);
csa_1509 csau_1509_i1322(tree_5[60359:58851],tree_5[61868:60360],tree_5[63377:61869],tree_6[40742:39234],tree_6[42251:40743]);
csa_1509 csau_1509_i1323(tree_5[64886:63378],tree_5[66395:64887],tree_5[67904:66396],tree_6[43760:42252],tree_6[45269:43761]);
csa_1509 csau_1509_i1324(tree_5[69413:67905],tree_5[70922:69414],tree_5[72431:70923],tree_6[46778:45270],tree_6[48287:46779]);
csa_1509 csau_1509_i1325(tree_5[73940:72432],tree_5[75449:73941],tree_5[76958:75450],tree_6[49796:48288],tree_6[51305:49797]);
csa_1509 csau_1509_i1326(tree_5[78467:76959],tree_5[79976:78468],tree_5[81485:79977],tree_6[52814:51306],tree_6[54323:52815]);
csa_1509 csau_1509_i1327(tree_5[82994:81486],tree_5[84503:82995],tree_5[86012:84504],tree_6[55832:54324],tree_6[57341:55833]);
csa_1509 csau_1509_i1328(tree_5[87521:86013],tree_5[89030:87522],tree_5[90539:89031],tree_6[58850:57342],tree_6[60359:58851]);
csa_1509 csau_1509_i1329(tree_5[92048:90540],tree_5[93557:92049],tree_5[95066:93558],tree_6[61868:60360],tree_6[63377:61869]);
csa_1509 csau_1509_i1330(tree_5[96575:95067],tree_5[98084:96576],tree_5[99593:98085],tree_6[64886:63378],tree_6[66395:64887]);
csa_1509 csau_1509_i1331(tree_5[101102:99594],tree_5[102611:101103],tree_5[104120:102612],tree_6[67904:66396],tree_6[69413:67905]);
csa_1509 csau_1509_i1332(tree_5[105629:104121],tree_5[107138:105630],tree_5[108647:107139],tree_6[70922:69414],tree_6[72431:70923]);
csa_1509 csau_1509_i1333(tree_5[110156:108648],tree_5[111665:110157],tree_5[113174:111666],tree_6[73940:72432],tree_6[75449:73941]);
csa_1509 csau_1509_i1334(tree_5[114683:113175],tree_5[116192:114684],tree_5[117701:116193],tree_6[76958:75450],tree_6[78467:76959]);
csa_1509 csau_1509_i1335(tree_5[119210:117702],tree_5[120719:119211],tree_5[122228:120720],tree_6[79976:78468],tree_6[81485:79977]);
csa_1509 csau_1509_i1336(tree_5[123737:122229],tree_5[125246:123738],tree_5[126755:125247],tree_6[82994:81486],tree_6[84503:82995]);
csa_1509 csau_1509_i1337(tree_5[128264:126756],tree_5[129773:128265],tree_5[131282:129774],tree_6[86012:84504],tree_6[87521:86013]);
csa_1509 csau_1509_i1338(tree_5[132791:131283],tree_5[134300:132792],tree_5[135809:134301],tree_6[89030:87522],tree_6[90539:89031]);
csa_1509 csau_1509_i1339(tree_5[137318:135810],tree_5[138827:137319],tree_5[140336:138828],tree_6[92048:90540],tree_6[93557:92049]);
csa_1509 csau_1509_i1340(tree_5[141845:140337],tree_5[143354:141846],tree_5[144863:143355],tree_6[95066:93558],tree_6[96575:95067]);
csa_1509 csau_1509_i1341(tree_5[146372:144864],tree_5[147881:146373],tree_5[149390:147882],tree_6[98084:96576],tree_6[99593:98085]);
csa_1509 csau_1509_i1342(tree_5[150899:149391],tree_5[152408:150900],tree_5[153917:152409],tree_6[101102:99594],tree_6[102611:101103]);
csa_1509 csau_1509_i1343(tree_5[155426:153918],tree_5[156935:155427],tree_5[158444:156936],tree_6[104120:102612],tree_6[105629:104121]);
csa_1509 csau_1509_i1344(tree_5[159953:158445],tree_5[161462:159954],tree_5[162971:161463],tree_6[107138:105630],tree_6[108647:107139]);
csa_1509 csau_1509_i1345(tree_5[164480:162972],tree_5[165989:164481],tree_5[167498:165990],tree_6[110156:108648],tree_6[111665:110157]);
csa_1509 csau_1509_i1346(tree_5[169007:167499],tree_5[170516:169008],tree_5[172025:170517],tree_6[113174:111666],tree_6[114683:113175]);
csa_1509 csau_1509_i1347(tree_5[173534:172026],tree_5[175043:173535],tree_5[176552:175044],tree_6[116192:114684],tree_6[117701:116193]);
csa_1509 csau_1509_i1348(tree_5[178061:176553],tree_5[179570:178062],tree_5[181079:179571],tree_6[119210:117702],tree_6[120719:119211]);
csa_1509 csau_1509_i1349(tree_5[182588:181080],tree_5[184097:182589],tree_5[185606:184098],tree_6[122228:120720],tree_6[123737:122229]);
csa_1509 csau_1509_i1350(tree_5[187115:185607],tree_5[188624:187116],tree_5[190133:188625],tree_6[125246:123738],tree_6[126755:125247]);
csa_1509 csau_1509_i1351(tree_5[191642:190134],tree_5[193151:191643],tree_5[194660:193152],tree_6[128264:126756],tree_6[129773:128265]);
csa_1509 csau_1509_i1352(tree_5[196169:194661],tree_5[197678:196170],tree_5[199187:197679],tree_6[131282:129774],tree_6[132791:131283]);
csa_1509 csau_1509_i1353(tree_5[200696:199188],tree_5[202205:200697],tree_5[203714:202206],tree_6[134300:132792],tree_6[135809:134301]);
csa_1509 csau_1509_i1354(tree_5[205223:203715],tree_5[206732:205224],tree_5[208241:206733],tree_6[137318:135810],tree_6[138827:137319]);
csa_1509 csau_1509_i1355(tree_5[209750:208242],tree_5[211259:209751],tree_5[212768:211260],tree_6[140336:138828],tree_6[141845:140337]);
csa_1509 csau_1509_i1356(tree_5[214277:212769],tree_5[215786:214278],tree_5[217295:215787],tree_6[143354:141846],tree_6[144863:143355]);
csa_1509 csau_1509_i1357(tree_5[218804:217296],tree_5[220313:218805],tree_5[221822:220314],tree_6[146372:144864],tree_6[147881:146373]);
csa_1509 csau_1509_i1358(tree_5[223331:221823],tree_5[224840:223332],tree_5[226349:224841],tree_6[149390:147882],tree_6[150899:149391]);
csa_1509 csau_1509_i1359(tree_5[227858:226350],tree_5[229367:227859],tree_5[230876:229368],tree_6[152408:150900],tree_6[153917:152409]);
csa_1509 csau_1509_i1360(tree_5[232385:230877],tree_5[233894:232386],tree_5[235403:233895],tree_6[155426:153918],tree_6[156935:155427]);
csa_1509 csau_1509_i1361(tree_5[236912:235404],tree_5[238421:236913],tree_5[239930:238422],tree_6[158444:156936],tree_6[159953:158445]);
csa_1509 csau_1509_i1362(tree_5[241439:239931],tree_5[242948:241440],tree_5[244457:242949],tree_6[161462:159954],tree_6[162971:161463]);
csa_1509 csau_1509_i1363(tree_5[245966:244458],tree_5[247475:245967],tree_5[248984:247476],tree_6[164480:162972],tree_6[165989:164481]);
csa_1509 csau_1509_i1364(tree_5[250493:248985],tree_5[252002:250494],tree_5[253511:252003],tree_6[167498:165990],tree_6[169007:167499]);
csa_1509 csau_1509_i1365(tree_5[255020:253512],tree_5[256529:255021],tree_5[258038:256530],tree_6[170516:169008],tree_6[172025:170517]);
csa_1509 csau_1509_i1366(tree_5[259547:258039],tree_5[261056:259548],tree_5[262565:261057],tree_6[173534:172026],tree_6[175043:173535]);
csa_1509 csau_1509_i1367(tree_5[264074:262566],tree_5[265583:264075],tree_5[267092:265584],tree_6[176552:175044],tree_6[178061:176553]);
csa_1509 csau_1509_i1368(tree_5[268601:267093],tree_5[270110:268602],tree_5[271619:270111],tree_6[179570:178062],tree_6[181079:179571]);
csa_1509 csau_1509_i1369(tree_5[273128:271620],tree_5[274637:273129],tree_5[276146:274638],tree_6[182588:181080],tree_6[184097:182589]);
csa_1509 csau_1509_i1370(tree_5[277655:276147],tree_5[279164:277656],tree_5[280673:279165],tree_6[185606:184098],tree_6[187115:185607]);
csa_1509 csau_1509_i1371(tree_5[282182:280674],tree_5[283691:282183],tree_5[285200:283692],tree_6[188624:187116],tree_6[190133:188625]);
csa_1509 csau_1509_i1372(tree_5[286709:285201],tree_5[288218:286710],tree_5[289727:288219],tree_6[191642:190134],tree_6[193151:191643]);
csa_1509 csau_1509_i1373(tree_5[291236:289728],tree_5[292745:291237],tree_5[294254:292746],tree_6[194660:193152],tree_6[196169:194661]);
csa_1509 csau_1509_i1374(tree_5[295763:294255],tree_5[297272:295764],tree_5[298781:297273],tree_6[197678:196170],tree_6[199187:197679]);
assign tree_6[200696:199188] = tree_5[300290:298782];
assign tree_6[202205:200697] = tree_5[301799:300291];
// layer-7
csa_1509 csau_1509_i1375(tree_6[1508:0],tree_6[3017:1509],tree_6[4526:3018],tree_7[1508:0],tree_7[3017:1509]);
csa_1509 csau_1509_i1376(tree_6[6035:4527],tree_6[7544:6036],tree_6[9053:7545],tree_7[4526:3018],tree_7[6035:4527]);
csa_1509 csau_1509_i1377(tree_6[10562:9054],tree_6[12071:10563],tree_6[13580:12072],tree_7[7544:6036],tree_7[9053:7545]);
csa_1509 csau_1509_i1378(tree_6[15089:13581],tree_6[16598:15090],tree_6[18107:16599],tree_7[10562:9054],tree_7[12071:10563]);
csa_1509 csau_1509_i1379(tree_6[19616:18108],tree_6[21125:19617],tree_6[22634:21126],tree_7[13580:12072],tree_7[15089:13581]);
csa_1509 csau_1509_i1380(tree_6[24143:22635],tree_6[25652:24144],tree_6[27161:25653],tree_7[16598:15090],tree_7[18107:16599]);
csa_1509 csau_1509_i1381(tree_6[28670:27162],tree_6[30179:28671],tree_6[31688:30180],tree_7[19616:18108],tree_7[21125:19617]);
csa_1509 csau_1509_i1382(tree_6[33197:31689],tree_6[34706:33198],tree_6[36215:34707],tree_7[22634:21126],tree_7[24143:22635]);
csa_1509 csau_1509_i1383(tree_6[37724:36216],tree_6[39233:37725],tree_6[40742:39234],tree_7[25652:24144],tree_7[27161:25653]);
csa_1509 csau_1509_i1384(tree_6[42251:40743],tree_6[43760:42252],tree_6[45269:43761],tree_7[28670:27162],tree_7[30179:28671]);
csa_1509 csau_1509_i1385(tree_6[46778:45270],tree_6[48287:46779],tree_6[49796:48288],tree_7[31688:30180],tree_7[33197:31689]);
csa_1509 csau_1509_i1386(tree_6[51305:49797],tree_6[52814:51306],tree_6[54323:52815],tree_7[34706:33198],tree_7[36215:34707]);
csa_1509 csau_1509_i1387(tree_6[55832:54324],tree_6[57341:55833],tree_6[58850:57342],tree_7[37724:36216],tree_7[39233:37725]);
csa_1509 csau_1509_i1388(tree_6[60359:58851],tree_6[61868:60360],tree_6[63377:61869],tree_7[40742:39234],tree_7[42251:40743]);
csa_1509 csau_1509_i1389(tree_6[64886:63378],tree_6[66395:64887],tree_6[67904:66396],tree_7[43760:42252],tree_7[45269:43761]);
csa_1509 csau_1509_i1390(tree_6[69413:67905],tree_6[70922:69414],tree_6[72431:70923],tree_7[46778:45270],tree_7[48287:46779]);
csa_1509 csau_1509_i1391(tree_6[73940:72432],tree_6[75449:73941],tree_6[76958:75450],tree_7[49796:48288],tree_7[51305:49797]);
csa_1509 csau_1509_i1392(tree_6[78467:76959],tree_6[79976:78468],tree_6[81485:79977],tree_7[52814:51306],tree_7[54323:52815]);
csa_1509 csau_1509_i1393(tree_6[82994:81486],tree_6[84503:82995],tree_6[86012:84504],tree_7[55832:54324],tree_7[57341:55833]);
csa_1509 csau_1509_i1394(tree_6[87521:86013],tree_6[89030:87522],tree_6[90539:89031],tree_7[58850:57342],tree_7[60359:58851]);
csa_1509 csau_1509_i1395(tree_6[92048:90540],tree_6[93557:92049],tree_6[95066:93558],tree_7[61868:60360],tree_7[63377:61869]);
csa_1509 csau_1509_i1396(tree_6[96575:95067],tree_6[98084:96576],tree_6[99593:98085],tree_7[64886:63378],tree_7[66395:64887]);
csa_1509 csau_1509_i1397(tree_6[101102:99594],tree_6[102611:101103],tree_6[104120:102612],tree_7[67904:66396],tree_7[69413:67905]);
csa_1509 csau_1509_i1398(tree_6[105629:104121],tree_6[107138:105630],tree_6[108647:107139],tree_7[70922:69414],tree_7[72431:70923]);
csa_1509 csau_1509_i1399(tree_6[110156:108648],tree_6[111665:110157],tree_6[113174:111666],tree_7[73940:72432],tree_7[75449:73941]);
csa_1509 csau_1509_i1400(tree_6[114683:113175],tree_6[116192:114684],tree_6[117701:116193],tree_7[76958:75450],tree_7[78467:76959]);
csa_1509 csau_1509_i1401(tree_6[119210:117702],tree_6[120719:119211],tree_6[122228:120720],tree_7[79976:78468],tree_7[81485:79977]);
csa_1509 csau_1509_i1402(tree_6[123737:122229],tree_6[125246:123738],tree_6[126755:125247],tree_7[82994:81486],tree_7[84503:82995]);
csa_1509 csau_1509_i1403(tree_6[128264:126756],tree_6[129773:128265],tree_6[131282:129774],tree_7[86012:84504],tree_7[87521:86013]);
csa_1509 csau_1509_i1404(tree_6[132791:131283],tree_6[134300:132792],tree_6[135809:134301],tree_7[89030:87522],tree_7[90539:89031]);
csa_1509 csau_1509_i1405(tree_6[137318:135810],tree_6[138827:137319],tree_6[140336:138828],tree_7[92048:90540],tree_7[93557:92049]);
csa_1509 csau_1509_i1406(tree_6[141845:140337],tree_6[143354:141846],tree_6[144863:143355],tree_7[95066:93558],tree_7[96575:95067]);
csa_1509 csau_1509_i1407(tree_6[146372:144864],tree_6[147881:146373],tree_6[149390:147882],tree_7[98084:96576],tree_7[99593:98085]);
csa_1509 csau_1509_i1408(tree_6[150899:149391],tree_6[152408:150900],tree_6[153917:152409],tree_7[101102:99594],tree_7[102611:101103]);
csa_1509 csau_1509_i1409(tree_6[155426:153918],tree_6[156935:155427],tree_6[158444:156936],tree_7[104120:102612],tree_7[105629:104121]);
csa_1509 csau_1509_i1410(tree_6[159953:158445],tree_6[161462:159954],tree_6[162971:161463],tree_7[107138:105630],tree_7[108647:107139]);
csa_1509 csau_1509_i1411(tree_6[164480:162972],tree_6[165989:164481],tree_6[167498:165990],tree_7[110156:108648],tree_7[111665:110157]);
csa_1509 csau_1509_i1412(tree_6[169007:167499],tree_6[170516:169008],tree_6[172025:170517],tree_7[113174:111666],tree_7[114683:113175]);
csa_1509 csau_1509_i1413(tree_6[173534:172026],tree_6[175043:173535],tree_6[176552:175044],tree_7[116192:114684],tree_7[117701:116193]);
csa_1509 csau_1509_i1414(tree_6[178061:176553],tree_6[179570:178062],tree_6[181079:179571],tree_7[119210:117702],tree_7[120719:119211]);
csa_1509 csau_1509_i1415(tree_6[182588:181080],tree_6[184097:182589],tree_6[185606:184098],tree_7[122228:120720],tree_7[123737:122229]);
csa_1509 csau_1509_i1416(tree_6[187115:185607],tree_6[188624:187116],tree_6[190133:188625],tree_7[125246:123738],tree_7[126755:125247]);
csa_1509 csau_1509_i1417(tree_6[191642:190134],tree_6[193151:191643],tree_6[194660:193152],tree_7[128264:126756],tree_7[129773:128265]);
csa_1509 csau_1509_i1418(tree_6[196169:194661],tree_6[197678:196170],tree_6[199187:197679],tree_7[131282:129774],tree_7[132791:131283]);
assign tree_7[134300:132792] = tree_6[200696:199188];
assign tree_7[135809:134301] = tree_6[202205:200697];
// layer-8
csa_1509 csau_1509_i1419(tree_7[1508:0],tree_7[3017:1509],tree_7[4526:3018],tree_8[1508:0],tree_8[3017:1509]);
csa_1509 csau_1509_i1420(tree_7[6035:4527],tree_7[7544:6036],tree_7[9053:7545],tree_8[4526:3018],tree_8[6035:4527]);
csa_1509 csau_1509_i1421(tree_7[10562:9054],tree_7[12071:10563],tree_7[13580:12072],tree_8[7544:6036],tree_8[9053:7545]);
csa_1509 csau_1509_i1422(tree_7[15089:13581],tree_7[16598:15090],tree_7[18107:16599],tree_8[10562:9054],tree_8[12071:10563]);
csa_1509 csau_1509_i1423(tree_7[19616:18108],tree_7[21125:19617],tree_7[22634:21126],tree_8[13580:12072],tree_8[15089:13581]);
csa_1509 csau_1509_i1424(tree_7[24143:22635],tree_7[25652:24144],tree_7[27161:25653],tree_8[16598:15090],tree_8[18107:16599]);
csa_1509 csau_1509_i1425(tree_7[28670:27162],tree_7[30179:28671],tree_7[31688:30180],tree_8[19616:18108],tree_8[21125:19617]);
csa_1509 csau_1509_i1426(tree_7[33197:31689],tree_7[34706:33198],tree_7[36215:34707],tree_8[22634:21126],tree_8[24143:22635]);
csa_1509 csau_1509_i1427(tree_7[37724:36216],tree_7[39233:37725],tree_7[40742:39234],tree_8[25652:24144],tree_8[27161:25653]);
csa_1509 csau_1509_i1428(tree_7[42251:40743],tree_7[43760:42252],tree_7[45269:43761],tree_8[28670:27162],tree_8[30179:28671]);
csa_1509 csau_1509_i1429(tree_7[46778:45270],tree_7[48287:46779],tree_7[49796:48288],tree_8[31688:30180],tree_8[33197:31689]);
csa_1509 csau_1509_i1430(tree_7[51305:49797],tree_7[52814:51306],tree_7[54323:52815],tree_8[34706:33198],tree_8[36215:34707]);
csa_1509 csau_1509_i1431(tree_7[55832:54324],tree_7[57341:55833],tree_7[58850:57342],tree_8[37724:36216],tree_8[39233:37725]);
csa_1509 csau_1509_i1432(tree_7[60359:58851],tree_7[61868:60360],tree_7[63377:61869],tree_8[40742:39234],tree_8[42251:40743]);
csa_1509 csau_1509_i1433(tree_7[64886:63378],tree_7[66395:64887],tree_7[67904:66396],tree_8[43760:42252],tree_8[45269:43761]);
csa_1509 csau_1509_i1434(tree_7[69413:67905],tree_7[70922:69414],tree_7[72431:70923],tree_8[46778:45270],tree_8[48287:46779]);
csa_1509 csau_1509_i1435(tree_7[73940:72432],tree_7[75449:73941],tree_7[76958:75450],tree_8[49796:48288],tree_8[51305:49797]);
csa_1509 csau_1509_i1436(tree_7[78467:76959],tree_7[79976:78468],tree_7[81485:79977],tree_8[52814:51306],tree_8[54323:52815]);
csa_1509 csau_1509_i1437(tree_7[82994:81486],tree_7[84503:82995],tree_7[86012:84504],tree_8[55832:54324],tree_8[57341:55833]);
csa_1509 csau_1509_i1438(tree_7[87521:86013],tree_7[89030:87522],tree_7[90539:89031],tree_8[58850:57342],tree_8[60359:58851]);
csa_1509 csau_1509_i1439(tree_7[92048:90540],tree_7[93557:92049],tree_7[95066:93558],tree_8[61868:60360],tree_8[63377:61869]);
csa_1509 csau_1509_i1440(tree_7[96575:95067],tree_7[98084:96576],tree_7[99593:98085],tree_8[64886:63378],tree_8[66395:64887]);
csa_1509 csau_1509_i1441(tree_7[101102:99594],tree_7[102611:101103],tree_7[104120:102612],tree_8[67904:66396],tree_8[69413:67905]);
csa_1509 csau_1509_i1442(tree_7[105629:104121],tree_7[107138:105630],tree_7[108647:107139],tree_8[70922:69414],tree_8[72431:70923]);
csa_1509 csau_1509_i1443(tree_7[110156:108648],tree_7[111665:110157],tree_7[113174:111666],tree_8[73940:72432],tree_8[75449:73941]);
csa_1509 csau_1509_i1444(tree_7[114683:113175],tree_7[116192:114684],tree_7[117701:116193],tree_8[76958:75450],tree_8[78467:76959]);
csa_1509 csau_1509_i1445(tree_7[119210:117702],tree_7[120719:119211],tree_7[122228:120720],tree_8[79976:78468],tree_8[81485:79977]);
csa_1509 csau_1509_i1446(tree_7[123737:122229],tree_7[125246:123738],tree_7[126755:125247],tree_8[82994:81486],tree_8[84503:82995]);
csa_1509 csau_1509_i1447(tree_7[128264:126756],tree_7[129773:128265],tree_7[131282:129774],tree_8[86012:84504],tree_8[87521:86013]);
csa_1509 csau_1509_i1448(tree_7[132791:131283],tree_7[134300:132792],tree_7[135809:134301],tree_8[89030:87522],tree_8[90539:89031]);
// layer-9
csa_1509 csau_1509_i1449(tree_8[1508:0],tree_8[3017:1509],tree_8[4526:3018],tree_9[1508:0],tree_9[3017:1509]);
csa_1509 csau_1509_i1450(tree_8[6035:4527],tree_8[7544:6036],tree_8[9053:7545],tree_9[4526:3018],tree_9[6035:4527]);
csa_1509 csau_1509_i1451(tree_8[10562:9054],tree_8[12071:10563],tree_8[13580:12072],tree_9[7544:6036],tree_9[9053:7545]);
csa_1509 csau_1509_i1452(tree_8[15089:13581],tree_8[16598:15090],tree_8[18107:16599],tree_9[10562:9054],tree_9[12071:10563]);
csa_1509 csau_1509_i1453(tree_8[19616:18108],tree_8[21125:19617],tree_8[22634:21126],tree_9[13580:12072],tree_9[15089:13581]);
csa_1509 csau_1509_i1454(tree_8[24143:22635],tree_8[25652:24144],tree_8[27161:25653],tree_9[16598:15090],tree_9[18107:16599]);
csa_1509 csau_1509_i1455(tree_8[28670:27162],tree_8[30179:28671],tree_8[31688:30180],tree_9[19616:18108],tree_9[21125:19617]);
csa_1509 csau_1509_i1456(tree_8[33197:31689],tree_8[34706:33198],tree_8[36215:34707],tree_9[22634:21126],tree_9[24143:22635]);
csa_1509 csau_1509_i1457(tree_8[37724:36216],tree_8[39233:37725],tree_8[40742:39234],tree_9[25652:24144],tree_9[27161:25653]);
csa_1509 csau_1509_i1458(tree_8[42251:40743],tree_8[43760:42252],tree_8[45269:43761],tree_9[28670:27162],tree_9[30179:28671]);
csa_1509 csau_1509_i1459(tree_8[46778:45270],tree_8[48287:46779],tree_8[49796:48288],tree_9[31688:30180],tree_9[33197:31689]);
csa_1509 csau_1509_i1460(tree_8[51305:49797],tree_8[52814:51306],tree_8[54323:52815],tree_9[34706:33198],tree_9[36215:34707]);
csa_1509 csau_1509_i1461(tree_8[55832:54324],tree_8[57341:55833],tree_8[58850:57342],tree_9[37724:36216],tree_9[39233:37725]);
csa_1509 csau_1509_i1462(tree_8[60359:58851],tree_8[61868:60360],tree_8[63377:61869],tree_9[40742:39234],tree_9[42251:40743]);
csa_1509 csau_1509_i1463(tree_8[64886:63378],tree_8[66395:64887],tree_8[67904:66396],tree_9[43760:42252],tree_9[45269:43761]);
csa_1509 csau_1509_i1464(tree_8[69413:67905],tree_8[70922:69414],tree_8[72431:70923],tree_9[46778:45270],tree_9[48287:46779]);
csa_1509 csau_1509_i1465(tree_8[73940:72432],tree_8[75449:73941],tree_8[76958:75450],tree_9[49796:48288],tree_9[51305:49797]);
csa_1509 csau_1509_i1466(tree_8[78467:76959],tree_8[79976:78468],tree_8[81485:79977],tree_9[52814:51306],tree_9[54323:52815]);
csa_1509 csau_1509_i1467(tree_8[82994:81486],tree_8[84503:82995],tree_8[86012:84504],tree_9[55832:54324],tree_9[57341:55833]);
csa_1509 csau_1509_i1468(tree_8[87521:86013],tree_8[89030:87522],tree_8[90539:89031],tree_9[58850:57342],tree_9[60359:58851]);
// layer-10
csa_1509 csau_1509_i1469(tree_9[1508:0],tree_9[3017:1509],tree_9[4526:3018],tree_10[1508:0],tree_10[3017:1509]);
csa_1509 csau_1509_i1470(tree_9[6035:4527],tree_9[7544:6036],tree_9[9053:7545],tree_10[4526:3018],tree_10[6035:4527]);
csa_1509 csau_1509_i1471(tree_9[10562:9054],tree_9[12071:10563],tree_9[13580:12072],tree_10[7544:6036],tree_10[9053:7545]);
csa_1509 csau_1509_i1472(tree_9[15089:13581],tree_9[16598:15090],tree_9[18107:16599],tree_10[10562:9054],tree_10[12071:10563]);
csa_1509 csau_1509_i1473(tree_9[19616:18108],tree_9[21125:19617],tree_9[22634:21126],tree_10[13580:12072],tree_10[15089:13581]);
csa_1509 csau_1509_i1474(tree_9[24143:22635],tree_9[25652:24144],tree_9[27161:25653],tree_10[16598:15090],tree_10[18107:16599]);
csa_1509 csau_1509_i1475(tree_9[28670:27162],tree_9[30179:28671],tree_9[31688:30180],tree_10[19616:18108],tree_10[21125:19617]);
csa_1509 csau_1509_i1476(tree_9[33197:31689],tree_9[34706:33198],tree_9[36215:34707],tree_10[22634:21126],tree_10[24143:22635]);
csa_1509 csau_1509_i1477(tree_9[37724:36216],tree_9[39233:37725],tree_9[40742:39234],tree_10[25652:24144],tree_10[27161:25653]);
csa_1509 csau_1509_i1478(tree_9[42251:40743],tree_9[43760:42252],tree_9[45269:43761],tree_10[28670:27162],tree_10[30179:28671]);
csa_1509 csau_1509_i1479(tree_9[46778:45270],tree_9[48287:46779],tree_9[49796:48288],tree_10[31688:30180],tree_10[33197:31689]);
csa_1509 csau_1509_i1480(tree_9[51305:49797],tree_9[52814:51306],tree_9[54323:52815],tree_10[34706:33198],tree_10[36215:34707]);
csa_1509 csau_1509_i1481(tree_9[55832:54324],tree_9[57341:55833],tree_9[58850:57342],tree_10[37724:36216],tree_10[39233:37725]);
assign tree_10[40742:39234] = tree_9[60359:58851];
// layer-11
csa_1509 csau_1509_i1482(tree_10[1508:0],tree_10[3017:1509],tree_10[4526:3018],tree_11[1508:0],tree_11[3017:1509]);
csa_1509 csau_1509_i1483(tree_10[6035:4527],tree_10[7544:6036],tree_10[9053:7545],tree_11[4526:3018],tree_11[6035:4527]);
csa_1509 csau_1509_i1484(tree_10[10562:9054],tree_10[12071:10563],tree_10[13580:12072],tree_11[7544:6036],tree_11[9053:7545]);
csa_1509 csau_1509_i1485(tree_10[15089:13581],tree_10[16598:15090],tree_10[18107:16599],tree_11[10562:9054],tree_11[12071:10563]);
csa_1509 csau_1509_i1486(tree_10[19616:18108],tree_10[21125:19617],tree_10[22634:21126],tree_11[13580:12072],tree_11[15089:13581]);
csa_1509 csau_1509_i1487(tree_10[24143:22635],tree_10[25652:24144],tree_10[27161:25653],tree_11[16598:15090],tree_11[18107:16599]);
csa_1509 csau_1509_i1488(tree_10[28670:27162],tree_10[30179:28671],tree_10[31688:30180],tree_11[19616:18108],tree_11[21125:19617]);
csa_1509 csau_1509_i1489(tree_10[33197:31689],tree_10[34706:33198],tree_10[36215:34707],tree_11[22634:21126],tree_11[24143:22635]);
csa_1509 csau_1509_i1490(tree_10[37724:36216],tree_10[39233:37725],tree_10[40742:39234],tree_11[25652:24144],tree_11[27161:25653]);
// layer-12
csa_1509 csau_1509_i1491(tree_11[1508:0],tree_11[3017:1509],tree_11[4526:3018],tree_12[1508:0],tree_12[3017:1509]);
csa_1509 csau_1509_i1492(tree_11[6035:4527],tree_11[7544:6036],tree_11[9053:7545],tree_12[4526:3018],tree_12[6035:4527]);
csa_1509 csau_1509_i1493(tree_11[10562:9054],tree_11[12071:10563],tree_11[13580:12072],tree_12[7544:6036],tree_12[9053:7545]);
csa_1509 csau_1509_i1494(tree_11[15089:13581],tree_11[16598:15090],tree_11[18107:16599],tree_12[10562:9054],tree_12[12071:10563]);
csa_1509 csau_1509_i1495(tree_11[19616:18108],tree_11[21125:19617],tree_11[22634:21126],tree_12[13580:12072],tree_12[15089:13581]);
csa_1509 csau_1509_i1496(tree_11[24143:22635],tree_11[25652:24144],tree_11[27161:25653],tree_12[16598:15090],tree_12[18107:16599]);
// layer-13
csa_1509 csau_1509_i1497(tree_12[1508:0],tree_12[3017:1509],tree_12[4526:3018],tree_13[1508:0],tree_13[3017:1509]);
csa_1509 csau_1509_i1498(tree_12[6035:4527],tree_12[7544:6036],tree_12[9053:7545],tree_13[4526:3018],tree_13[6035:4527]);
csa_1509 csau_1509_i1499(tree_12[10562:9054],tree_12[12071:10563],tree_12[13580:12072],tree_13[7544:6036],tree_13[9053:7545]);
csa_1509 csau_1509_i1500(tree_12[15089:13581],tree_12[16598:15090],tree_12[18107:16599],tree_13[10562:9054],tree_13[12071:10563]);
// layer-14
csa_1509 csau_1509_i1501(tree_13[1508:0],tree_13[3017:1509],tree_13[4526:3018],tree_14[1508:0],tree_14[3017:1509]);
csa_1509 csau_1509_i1502(tree_13[6035:4527],tree_13[7544:6036],tree_13[9053:7545],tree_14[4526:3018],tree_14[6035:4527]);
assign tree_14[7544:6036] = tree_13[10562:9054];
assign tree_14[9053:7545] = tree_13[12071:10563];
// layer-15
csa_1509 csau_1509_i1503(tree_14[1508:0],tree_14[3017:1509],tree_14[4526:3018],tree_15[1508:0],tree_15[3017:1509]);
csa_1509 csau_1509_i1504(tree_14[6035:4527],tree_14[7544:6036],tree_14[9053:7545],tree_15[4526:3018],tree_15[6035:4527]);
// layer-16
csa_1509 csau_1509_i1505(tree_15[1508:0],tree_15[3017:1509],tree_15[4526:3018],tree_16[1508:0],tree_16[3017:1509]);
assign tree_16[4526:3018] = tree_15[6035:4527];
// layer-17
csa_1509 csau_1509_i1506(tree_16[1508:0],tree_16[3017:1509],tree_16[4526:3018],tree_17[1508:0],tree_17[3017:1509]);

// final assignment
assign B_0 = tree_17[1508:0];
assign B_1 = tree_17[3017:1509];

endmodule
