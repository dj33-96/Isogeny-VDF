
module red_part1_1509x1509(
    input [3013:0] a_c,a_s,
    input [1508:0] p_prime,
    output [2277080:0] b_c,b_s // lines are appended together
);
    
wire [1508:0] c_w_0, s_w_0;
wire [1508:0] c_w_1, s_w_1;
wire [1508:0] c_w_2, s_w_2;
wire [1508:0] c_w_3, s_w_3;
wire [1508:0] c_w_4, s_w_4;
wire [1508:0] c_w_5, s_w_5;
wire [1508:0] c_w_6, s_w_6;
wire [1508:0] c_w_7, s_w_7;
wire [1508:0] c_w_8, s_w_8;
wire [1508:0] c_w_9, s_w_9;
wire [1508:0] c_w_10, s_w_10;
wire [1508:0] c_w_11, s_w_11;
wire [1508:0] c_w_12, s_w_12;
wire [1508:0] c_w_13, s_w_13;
wire [1508:0] c_w_14, s_w_14;
wire [1508:0] c_w_15, s_w_15;
wire [1508:0] c_w_16, s_w_16;
wire [1508:0] c_w_17, s_w_17;
wire [1508:0] c_w_18, s_w_18;
wire [1508:0] c_w_19, s_w_19;
wire [1508:0] c_w_20, s_w_20;
wire [1508:0] c_w_21, s_w_21;
wire [1508:0] c_w_22, s_w_22;
wire [1508:0] c_w_23, s_w_23;
wire [1508:0] c_w_24, s_w_24;
wire [1508:0] c_w_25, s_w_25;
wire [1508:0] c_w_26, s_w_26;
wire [1508:0] c_w_27, s_w_27;
wire [1508:0] c_w_28, s_w_28;
wire [1508:0] c_w_29, s_w_29;
wire [1508:0] c_w_30, s_w_30;
wire [1508:0] c_w_31, s_w_31;
wire [1508:0] c_w_32, s_w_32;
wire [1508:0] c_w_33, s_w_33;
wire [1508:0] c_w_34, s_w_34;
wire [1508:0] c_w_35, s_w_35;
wire [1508:0] c_w_36, s_w_36;
wire [1508:0] c_w_37, s_w_37;
wire [1508:0] c_w_38, s_w_38;
wire [1508:0] c_w_39, s_w_39;
wire [1508:0] c_w_40, s_w_40;
wire [1508:0] c_w_41, s_w_41;
wire [1508:0] c_w_42, s_w_42;
wire [1508:0] c_w_43, s_w_43;
wire [1508:0] c_w_44, s_w_44;
wire [1508:0] c_w_45, s_w_45;
wire [1508:0] c_w_46, s_w_46;
wire [1508:0] c_w_47, s_w_47;
wire [1508:0] c_w_48, s_w_48;
wire [1508:0] c_w_49, s_w_49;
wire [1508:0] c_w_50, s_w_50;
wire [1508:0] c_w_51, s_w_51;
wire [1508:0] c_w_52, s_w_52;
wire [1508:0] c_w_53, s_w_53;
wire [1508:0] c_w_54, s_w_54;
wire [1508:0] c_w_55, s_w_55;
wire [1508:0] c_w_56, s_w_56;
wire [1508:0] c_w_57, s_w_57;
wire [1508:0] c_w_58, s_w_58;
wire [1508:0] c_w_59, s_w_59;
wire [1508:0] c_w_60, s_w_60;
wire [1508:0] c_w_61, s_w_61;
wire [1508:0] c_w_62, s_w_62;
wire [1508:0] c_w_63, s_w_63;
wire [1508:0] c_w_64, s_w_64;
wire [1508:0] c_w_65, s_w_65;
wire [1508:0] c_w_66, s_w_66;
wire [1508:0] c_w_67, s_w_67;
wire [1508:0] c_w_68, s_w_68;
wire [1508:0] c_w_69, s_w_69;
wire [1508:0] c_w_70, s_w_70;
wire [1508:0] c_w_71, s_w_71;
wire [1508:0] c_w_72, s_w_72;
wire [1508:0] c_w_73, s_w_73;
wire [1508:0] c_w_74, s_w_74;
wire [1508:0] c_w_75, s_w_75;
wire [1508:0] c_w_76, s_w_76;
wire [1508:0] c_w_77, s_w_77;
wire [1508:0] c_w_78, s_w_78;
wire [1508:0] c_w_79, s_w_79;
wire [1508:0] c_w_80, s_w_80;
wire [1508:0] c_w_81, s_w_81;
wire [1508:0] c_w_82, s_w_82;
wire [1508:0] c_w_83, s_w_83;
wire [1508:0] c_w_84, s_w_84;
wire [1508:0] c_w_85, s_w_85;
wire [1508:0] c_w_86, s_w_86;
wire [1508:0] c_w_87, s_w_87;
wire [1508:0] c_w_88, s_w_88;
wire [1508:0] c_w_89, s_w_89;
wire [1508:0] c_w_90, s_w_90;
wire [1508:0] c_w_91, s_w_91;
wire [1508:0] c_w_92, s_w_92;
wire [1508:0] c_w_93, s_w_93;
wire [1508:0] c_w_94, s_w_94;
wire [1508:0] c_w_95, s_w_95;
wire [1508:0] c_w_96, s_w_96;
wire [1508:0] c_w_97, s_w_97;
wire [1508:0] c_w_98, s_w_98;
wire [1508:0] c_w_99, s_w_99;
wire [1508:0] c_w_100, s_w_100;
wire [1508:0] c_w_101, s_w_101;
wire [1508:0] c_w_102, s_w_102;
wire [1508:0] c_w_103, s_w_103;
wire [1508:0] c_w_104, s_w_104;
wire [1508:0] c_w_105, s_w_105;
wire [1508:0] c_w_106, s_w_106;
wire [1508:0] c_w_107, s_w_107;
wire [1508:0] c_w_108, s_w_108;
wire [1508:0] c_w_109, s_w_109;
wire [1508:0] c_w_110, s_w_110;
wire [1508:0] c_w_111, s_w_111;
wire [1508:0] c_w_112, s_w_112;
wire [1508:0] c_w_113, s_w_113;
wire [1508:0] c_w_114, s_w_114;
wire [1508:0] c_w_115, s_w_115;
wire [1508:0] c_w_116, s_w_116;
wire [1508:0] c_w_117, s_w_117;
wire [1508:0] c_w_118, s_w_118;
wire [1508:0] c_w_119, s_w_119;
wire [1508:0] c_w_120, s_w_120;
wire [1508:0] c_w_121, s_w_121;
wire [1508:0] c_w_122, s_w_122;
wire [1508:0] c_w_123, s_w_123;
wire [1508:0] c_w_124, s_w_124;
wire [1508:0] c_w_125, s_w_125;
wire [1508:0] c_w_126, s_w_126;
wire [1508:0] c_w_127, s_w_127;
wire [1508:0] c_w_128, s_w_128;
wire [1508:0] c_w_129, s_w_129;
wire [1508:0] c_w_130, s_w_130;
wire [1508:0] c_w_131, s_w_131;
wire [1508:0] c_w_132, s_w_132;
wire [1508:0] c_w_133, s_w_133;
wire [1508:0] c_w_134, s_w_134;
wire [1508:0] c_w_135, s_w_135;
wire [1508:0] c_w_136, s_w_136;
wire [1508:0] c_w_137, s_w_137;
wire [1508:0] c_w_138, s_w_138;
wire [1508:0] c_w_139, s_w_139;
wire [1508:0] c_w_140, s_w_140;
wire [1508:0] c_w_141, s_w_141;
wire [1508:0] c_w_142, s_w_142;
wire [1508:0] c_w_143, s_w_143;
wire [1508:0] c_w_144, s_w_144;
wire [1508:0] c_w_145, s_w_145;
wire [1508:0] c_w_146, s_w_146;
wire [1508:0] c_w_147, s_w_147;
wire [1508:0] c_w_148, s_w_148;
wire [1508:0] c_w_149, s_w_149;
wire [1508:0] c_w_150, s_w_150;
wire [1508:0] c_w_151, s_w_151;
wire [1508:0] c_w_152, s_w_152;
wire [1508:0] c_w_153, s_w_153;
wire [1508:0] c_w_154, s_w_154;
wire [1508:0] c_w_155, s_w_155;
wire [1508:0] c_w_156, s_w_156;
wire [1508:0] c_w_157, s_w_157;
wire [1508:0] c_w_158, s_w_158;
wire [1508:0] c_w_159, s_w_159;
wire [1508:0] c_w_160, s_w_160;
wire [1508:0] c_w_161, s_w_161;
wire [1508:0] c_w_162, s_w_162;
wire [1508:0] c_w_163, s_w_163;
wire [1508:0] c_w_164, s_w_164;
wire [1508:0] c_w_165, s_w_165;
wire [1508:0] c_w_166, s_w_166;
wire [1508:0] c_w_167, s_w_167;
wire [1508:0] c_w_168, s_w_168;
wire [1508:0] c_w_169, s_w_169;
wire [1508:0] c_w_170, s_w_170;
wire [1508:0] c_w_171, s_w_171;
wire [1508:0] c_w_172, s_w_172;
wire [1508:0] c_w_173, s_w_173;
wire [1508:0] c_w_174, s_w_174;
wire [1508:0] c_w_175, s_w_175;
wire [1508:0] c_w_176, s_w_176;
wire [1508:0] c_w_177, s_w_177;
wire [1508:0] c_w_178, s_w_178;
wire [1508:0] c_w_179, s_w_179;
wire [1508:0] c_w_180, s_w_180;
wire [1508:0] c_w_181, s_w_181;
wire [1508:0] c_w_182, s_w_182;
wire [1508:0] c_w_183, s_w_183;
wire [1508:0] c_w_184, s_w_184;
wire [1508:0] c_w_185, s_w_185;
wire [1508:0] c_w_186, s_w_186;
wire [1508:0] c_w_187, s_w_187;
wire [1508:0] c_w_188, s_w_188;
wire [1508:0] c_w_189, s_w_189;
wire [1508:0] c_w_190, s_w_190;
wire [1508:0] c_w_191, s_w_191;
wire [1508:0] c_w_192, s_w_192;
wire [1508:0] c_w_193, s_w_193;
wire [1508:0] c_w_194, s_w_194;
wire [1508:0] c_w_195, s_w_195;
wire [1508:0] c_w_196, s_w_196;
wire [1508:0] c_w_197, s_w_197;
wire [1508:0] c_w_198, s_w_198;
wire [1508:0] c_w_199, s_w_199;
wire [1508:0] c_w_200, s_w_200;
wire [1508:0] c_w_201, s_w_201;
wire [1508:0] c_w_202, s_w_202;
wire [1508:0] c_w_203, s_w_203;
wire [1508:0] c_w_204, s_w_204;
wire [1508:0] c_w_205, s_w_205;
wire [1508:0] c_w_206, s_w_206;
wire [1508:0] c_w_207, s_w_207;
wire [1508:0] c_w_208, s_w_208;
wire [1508:0] c_w_209, s_w_209;
wire [1508:0] c_w_210, s_w_210;
wire [1508:0] c_w_211, s_w_211;
wire [1508:0] c_w_212, s_w_212;
wire [1508:0] c_w_213, s_w_213;
wire [1508:0] c_w_214, s_w_214;
wire [1508:0] c_w_215, s_w_215;
wire [1508:0] c_w_216, s_w_216;
wire [1508:0] c_w_217, s_w_217;
wire [1508:0] c_w_218, s_w_218;
wire [1508:0] c_w_219, s_w_219;
wire [1508:0] c_w_220, s_w_220;
wire [1508:0] c_w_221, s_w_221;
wire [1508:0] c_w_222, s_w_222;
wire [1508:0] c_w_223, s_w_223;
wire [1508:0] c_w_224, s_w_224;
wire [1508:0] c_w_225, s_w_225;
wire [1508:0] c_w_226, s_w_226;
wire [1508:0] c_w_227, s_w_227;
wire [1508:0] c_w_228, s_w_228;
wire [1508:0] c_w_229, s_w_229;
wire [1508:0] c_w_230, s_w_230;
wire [1508:0] c_w_231, s_w_231;
wire [1508:0] c_w_232, s_w_232;
wire [1508:0] c_w_233, s_w_233;
wire [1508:0] c_w_234, s_w_234;
wire [1508:0] c_w_235, s_w_235;
wire [1508:0] c_w_236, s_w_236;
wire [1508:0] c_w_237, s_w_237;
wire [1508:0] c_w_238, s_w_238;
wire [1508:0] c_w_239, s_w_239;
wire [1508:0] c_w_240, s_w_240;
wire [1508:0] c_w_241, s_w_241;
wire [1508:0] c_w_242, s_w_242;
wire [1508:0] c_w_243, s_w_243;
wire [1508:0] c_w_244, s_w_244;
wire [1508:0] c_w_245, s_w_245;
wire [1508:0] c_w_246, s_w_246;
wire [1508:0] c_w_247, s_w_247;
wire [1508:0] c_w_248, s_w_248;
wire [1508:0] c_w_249, s_w_249;
wire [1508:0] c_w_250, s_w_250;
wire [1508:0] c_w_251, s_w_251;
wire [1508:0] c_w_252, s_w_252;
wire [1508:0] c_w_253, s_w_253;
wire [1508:0] c_w_254, s_w_254;
wire [1508:0] c_w_255, s_w_255;
wire [1508:0] c_w_256, s_w_256;
wire [1508:0] c_w_257, s_w_257;
wire [1508:0] c_w_258, s_w_258;
wire [1508:0] c_w_259, s_w_259;
wire [1508:0] c_w_260, s_w_260;
wire [1508:0] c_w_261, s_w_261;
wire [1508:0] c_w_262, s_w_262;
wire [1508:0] c_w_263, s_w_263;
wire [1508:0] c_w_264, s_w_264;
wire [1508:0] c_w_265, s_w_265;
wire [1508:0] c_w_266, s_w_266;
wire [1508:0] c_w_267, s_w_267;
wire [1508:0] c_w_268, s_w_268;
wire [1508:0] c_w_269, s_w_269;
wire [1508:0] c_w_270, s_w_270;
wire [1508:0] c_w_271, s_w_271;
wire [1508:0] c_w_272, s_w_272;
wire [1508:0] c_w_273, s_w_273;
wire [1508:0] c_w_274, s_w_274;
wire [1508:0] c_w_275, s_w_275;
wire [1508:0] c_w_276, s_w_276;
wire [1508:0] c_w_277, s_w_277;
wire [1508:0] c_w_278, s_w_278;
wire [1508:0] c_w_279, s_w_279;
wire [1508:0] c_w_280, s_w_280;
wire [1508:0] c_w_281, s_w_281;
wire [1508:0] c_w_282, s_w_282;
wire [1508:0] c_w_283, s_w_283;
wire [1508:0] c_w_284, s_w_284;
wire [1508:0] c_w_285, s_w_285;
wire [1508:0] c_w_286, s_w_286;
wire [1508:0] c_w_287, s_w_287;
wire [1508:0] c_w_288, s_w_288;
wire [1508:0] c_w_289, s_w_289;
wire [1508:0] c_w_290, s_w_290;
wire [1508:0] c_w_291, s_w_291;
wire [1508:0] c_w_292, s_w_292;
wire [1508:0] c_w_293, s_w_293;
wire [1508:0] c_w_294, s_w_294;
wire [1508:0] c_w_295, s_w_295;
wire [1508:0] c_w_296, s_w_296;
wire [1508:0] c_w_297, s_w_297;
wire [1508:0] c_w_298, s_w_298;
wire [1508:0] c_w_299, s_w_299;
wire [1508:0] c_w_300, s_w_300;
wire [1508:0] c_w_301, s_w_301;
wire [1508:0] c_w_302, s_w_302;
wire [1508:0] c_w_303, s_w_303;
wire [1508:0] c_w_304, s_w_304;
wire [1508:0] c_w_305, s_w_305;
wire [1508:0] c_w_306, s_w_306;
wire [1508:0] c_w_307, s_w_307;
wire [1508:0] c_w_308, s_w_308;
wire [1508:0] c_w_309, s_w_309;
wire [1508:0] c_w_310, s_w_310;
wire [1508:0] c_w_311, s_w_311;
wire [1508:0] c_w_312, s_w_312;
wire [1508:0] c_w_313, s_w_313;
wire [1508:0] c_w_314, s_w_314;
wire [1508:0] c_w_315, s_w_315;
wire [1508:0] c_w_316, s_w_316;
wire [1508:0] c_w_317, s_w_317;
wire [1508:0] c_w_318, s_w_318;
wire [1508:0] c_w_319, s_w_319;
wire [1508:0] c_w_320, s_w_320;
wire [1508:0] c_w_321, s_w_321;
wire [1508:0] c_w_322, s_w_322;
wire [1508:0] c_w_323, s_w_323;
wire [1508:0] c_w_324, s_w_324;
wire [1508:0] c_w_325, s_w_325;
wire [1508:0] c_w_326, s_w_326;
wire [1508:0] c_w_327, s_w_327;
wire [1508:0] c_w_328, s_w_328;
wire [1508:0] c_w_329, s_w_329;
wire [1508:0] c_w_330, s_w_330;
wire [1508:0] c_w_331, s_w_331;
wire [1508:0] c_w_332, s_w_332;
wire [1508:0] c_w_333, s_w_333;
wire [1508:0] c_w_334, s_w_334;
wire [1508:0] c_w_335, s_w_335;
wire [1508:0] c_w_336, s_w_336;
wire [1508:0] c_w_337, s_w_337;
wire [1508:0] c_w_338, s_w_338;
wire [1508:0] c_w_339, s_w_339;
wire [1508:0] c_w_340, s_w_340;
wire [1508:0] c_w_341, s_w_341;
wire [1508:0] c_w_342, s_w_342;
wire [1508:0] c_w_343, s_w_343;
wire [1508:0] c_w_344, s_w_344;
wire [1508:0] c_w_345, s_w_345;
wire [1508:0] c_w_346, s_w_346;
wire [1508:0] c_w_347, s_w_347;
wire [1508:0] c_w_348, s_w_348;
wire [1508:0] c_w_349, s_w_349;
wire [1508:0] c_w_350, s_w_350;
wire [1508:0] c_w_351, s_w_351;
wire [1508:0] c_w_352, s_w_352;
wire [1508:0] c_w_353, s_w_353;
wire [1508:0] c_w_354, s_w_354;
wire [1508:0] c_w_355, s_w_355;
wire [1508:0] c_w_356, s_w_356;
wire [1508:0] c_w_357, s_w_357;
wire [1508:0] c_w_358, s_w_358;
wire [1508:0] c_w_359, s_w_359;
wire [1508:0] c_w_360, s_w_360;
wire [1508:0] c_w_361, s_w_361;
wire [1508:0] c_w_362, s_w_362;
wire [1508:0] c_w_363, s_w_363;
wire [1508:0] c_w_364, s_w_364;
wire [1508:0] c_w_365, s_w_365;
wire [1508:0] c_w_366, s_w_366;
wire [1508:0] c_w_367, s_w_367;
wire [1508:0] c_w_368, s_w_368;
wire [1508:0] c_w_369, s_w_369;
wire [1508:0] c_w_370, s_w_370;
wire [1508:0] c_w_371, s_w_371;
wire [1508:0] c_w_372, s_w_372;
wire [1508:0] c_w_373, s_w_373;
wire [1508:0] c_w_374, s_w_374;
wire [1508:0] c_w_375, s_w_375;
wire [1508:0] c_w_376, s_w_376;
wire [1508:0] c_w_377, s_w_377;
wire [1508:0] c_w_378, s_w_378;
wire [1508:0] c_w_379, s_w_379;
wire [1508:0] c_w_380, s_w_380;
wire [1508:0] c_w_381, s_w_381;
wire [1508:0] c_w_382, s_w_382;
wire [1508:0] c_w_383, s_w_383;
wire [1508:0] c_w_384, s_w_384;
wire [1508:0] c_w_385, s_w_385;
wire [1508:0] c_w_386, s_w_386;
wire [1508:0] c_w_387, s_w_387;
wire [1508:0] c_w_388, s_w_388;
wire [1508:0] c_w_389, s_w_389;
wire [1508:0] c_w_390, s_w_390;
wire [1508:0] c_w_391, s_w_391;
wire [1508:0] c_w_392, s_w_392;
wire [1508:0] c_w_393, s_w_393;
wire [1508:0] c_w_394, s_w_394;
wire [1508:0] c_w_395, s_w_395;
wire [1508:0] c_w_396, s_w_396;
wire [1508:0] c_w_397, s_w_397;
wire [1508:0] c_w_398, s_w_398;
wire [1508:0] c_w_399, s_w_399;
wire [1508:0] c_w_400, s_w_400;
wire [1508:0] c_w_401, s_w_401;
wire [1508:0] c_w_402, s_w_402;
wire [1508:0] c_w_403, s_w_403;
wire [1508:0] c_w_404, s_w_404;
wire [1508:0] c_w_405, s_w_405;
wire [1508:0] c_w_406, s_w_406;
wire [1508:0] c_w_407, s_w_407;
wire [1508:0] c_w_408, s_w_408;
wire [1508:0] c_w_409, s_w_409;
wire [1508:0] c_w_410, s_w_410;
wire [1508:0] c_w_411, s_w_411;
wire [1508:0] c_w_412, s_w_412;
wire [1508:0] c_w_413, s_w_413;
wire [1508:0] c_w_414, s_w_414;
wire [1508:0] c_w_415, s_w_415;
wire [1508:0] c_w_416, s_w_416;
wire [1508:0] c_w_417, s_w_417;
wire [1508:0] c_w_418, s_w_418;
wire [1508:0] c_w_419, s_w_419;
wire [1508:0] c_w_420, s_w_420;
wire [1508:0] c_w_421, s_w_421;
wire [1508:0] c_w_422, s_w_422;
wire [1508:0] c_w_423, s_w_423;
wire [1508:0] c_w_424, s_w_424;
wire [1508:0] c_w_425, s_w_425;
wire [1508:0] c_w_426, s_w_426;
wire [1508:0] c_w_427, s_w_427;
wire [1508:0] c_w_428, s_w_428;
wire [1508:0] c_w_429, s_w_429;
wire [1508:0] c_w_430, s_w_430;
wire [1508:0] c_w_431, s_w_431;
wire [1508:0] c_w_432, s_w_432;
wire [1508:0] c_w_433, s_w_433;
wire [1508:0] c_w_434, s_w_434;
wire [1508:0] c_w_435, s_w_435;
wire [1508:0] c_w_436, s_w_436;
wire [1508:0] c_w_437, s_w_437;
wire [1508:0] c_w_438, s_w_438;
wire [1508:0] c_w_439, s_w_439;
wire [1508:0] c_w_440, s_w_440;
wire [1508:0] c_w_441, s_w_441;
wire [1508:0] c_w_442, s_w_442;
wire [1508:0] c_w_443, s_w_443;
wire [1508:0] c_w_444, s_w_444;
wire [1508:0] c_w_445, s_w_445;
wire [1508:0] c_w_446, s_w_446;
wire [1508:0] c_w_447, s_w_447;
wire [1508:0] c_w_448, s_w_448;
wire [1508:0] c_w_449, s_w_449;
wire [1508:0] c_w_450, s_w_450;
wire [1508:0] c_w_451, s_w_451;
wire [1508:0] c_w_452, s_w_452;
wire [1508:0] c_w_453, s_w_453;
wire [1508:0] c_w_454, s_w_454;
wire [1508:0] c_w_455, s_w_455;
wire [1508:0] c_w_456, s_w_456;
wire [1508:0] c_w_457, s_w_457;
wire [1508:0] c_w_458, s_w_458;
wire [1508:0] c_w_459, s_w_459;
wire [1508:0] c_w_460, s_w_460;
wire [1508:0] c_w_461, s_w_461;
wire [1508:0] c_w_462, s_w_462;
wire [1508:0] c_w_463, s_w_463;
wire [1508:0] c_w_464, s_w_464;
wire [1508:0] c_w_465, s_w_465;
wire [1508:0] c_w_466, s_w_466;
wire [1508:0] c_w_467, s_w_467;
wire [1508:0] c_w_468, s_w_468;
wire [1508:0] c_w_469, s_w_469;
wire [1508:0] c_w_470, s_w_470;
wire [1508:0] c_w_471, s_w_471;
wire [1508:0] c_w_472, s_w_472;
wire [1508:0] c_w_473, s_w_473;
wire [1508:0] c_w_474, s_w_474;
wire [1508:0] c_w_475, s_w_475;
wire [1508:0] c_w_476, s_w_476;
wire [1508:0] c_w_477, s_w_477;
wire [1508:0] c_w_478, s_w_478;
wire [1508:0] c_w_479, s_w_479;
wire [1508:0] c_w_480, s_w_480;
wire [1508:0] c_w_481, s_w_481;
wire [1508:0] c_w_482, s_w_482;
wire [1508:0] c_w_483, s_w_483;
wire [1508:0] c_w_484, s_w_484;
wire [1508:0] c_w_485, s_w_485;
wire [1508:0] c_w_486, s_w_486;
wire [1508:0] c_w_487, s_w_487;
wire [1508:0] c_w_488, s_w_488;
wire [1508:0] c_w_489, s_w_489;
wire [1508:0] c_w_490, s_w_490;
wire [1508:0] c_w_491, s_w_491;
wire [1508:0] c_w_492, s_w_492;
wire [1508:0] c_w_493, s_w_493;
wire [1508:0] c_w_494, s_w_494;
wire [1508:0] c_w_495, s_w_495;
wire [1508:0] c_w_496, s_w_496;
wire [1508:0] c_w_497, s_w_497;
wire [1508:0] c_w_498, s_w_498;
wire [1508:0] c_w_499, s_w_499;
wire [1508:0] c_w_500, s_w_500;
wire [1508:0] c_w_501, s_w_501;
wire [1508:0] c_w_502, s_w_502;
wire [1508:0] c_w_503, s_w_503;
wire [1508:0] c_w_504, s_w_504;
wire [1508:0] c_w_505, s_w_505;
wire [1508:0] c_w_506, s_w_506;
wire [1508:0] c_w_507, s_w_507;
wire [1508:0] c_w_508, s_w_508;
wire [1508:0] c_w_509, s_w_509;
wire [1508:0] c_w_510, s_w_510;
wire [1508:0] c_w_511, s_w_511;
wire [1508:0] c_w_512, s_w_512;
wire [1508:0] c_w_513, s_w_513;
wire [1508:0] c_w_514, s_w_514;
wire [1508:0] c_w_515, s_w_515;
wire [1508:0] c_w_516, s_w_516;
wire [1508:0] c_w_517, s_w_517;
wire [1508:0] c_w_518, s_w_518;
wire [1508:0] c_w_519, s_w_519;
wire [1508:0] c_w_520, s_w_520;
wire [1508:0] c_w_521, s_w_521;
wire [1508:0] c_w_522, s_w_522;
wire [1508:0] c_w_523, s_w_523;
wire [1508:0] c_w_524, s_w_524;
wire [1508:0] c_w_525, s_w_525;
wire [1508:0] c_w_526, s_w_526;
wire [1508:0] c_w_527, s_w_527;
wire [1508:0] c_w_528, s_w_528;
wire [1508:0] c_w_529, s_w_529;
wire [1508:0] c_w_530, s_w_530;
wire [1508:0] c_w_531, s_w_531;
wire [1508:0] c_w_532, s_w_532;
wire [1508:0] c_w_533, s_w_533;
wire [1508:0] c_w_534, s_w_534;
wire [1508:0] c_w_535, s_w_535;
wire [1508:0] c_w_536, s_w_536;
wire [1508:0] c_w_537, s_w_537;
wire [1508:0] c_w_538, s_w_538;
wire [1508:0] c_w_539, s_w_539;
wire [1508:0] c_w_540, s_w_540;
wire [1508:0] c_w_541, s_w_541;
wire [1508:0] c_w_542, s_w_542;
wire [1508:0] c_w_543, s_w_543;
wire [1508:0] c_w_544, s_w_544;
wire [1508:0] c_w_545, s_w_545;
wire [1508:0] c_w_546, s_w_546;
wire [1508:0] c_w_547, s_w_547;
wire [1508:0] c_w_548, s_w_548;
wire [1508:0] c_w_549, s_w_549;
wire [1508:0] c_w_550, s_w_550;
wire [1508:0] c_w_551, s_w_551;
wire [1508:0] c_w_552, s_w_552;
wire [1508:0] c_w_553, s_w_553;
wire [1508:0] c_w_554, s_w_554;
wire [1508:0] c_w_555, s_w_555;
wire [1508:0] c_w_556, s_w_556;
wire [1508:0] c_w_557, s_w_557;
wire [1508:0] c_w_558, s_w_558;
wire [1508:0] c_w_559, s_w_559;
wire [1508:0] c_w_560, s_w_560;
wire [1508:0] c_w_561, s_w_561;
wire [1508:0] c_w_562, s_w_562;
wire [1508:0] c_w_563, s_w_563;
wire [1508:0] c_w_564, s_w_564;
wire [1508:0] c_w_565, s_w_565;
wire [1508:0] c_w_566, s_w_566;
wire [1508:0] c_w_567, s_w_567;
wire [1508:0] c_w_568, s_w_568;
wire [1508:0] c_w_569, s_w_569;
wire [1508:0] c_w_570, s_w_570;
wire [1508:0] c_w_571, s_w_571;
wire [1508:0] c_w_572, s_w_572;
wire [1508:0] c_w_573, s_w_573;
wire [1508:0] c_w_574, s_w_574;
wire [1508:0] c_w_575, s_w_575;
wire [1508:0] c_w_576, s_w_576;
wire [1508:0] c_w_577, s_w_577;
wire [1508:0] c_w_578, s_w_578;
wire [1508:0] c_w_579, s_w_579;
wire [1508:0] c_w_580, s_w_580;
wire [1508:0] c_w_581, s_w_581;
wire [1508:0] c_w_582, s_w_582;
wire [1508:0] c_w_583, s_w_583;
wire [1508:0] c_w_584, s_w_584;
wire [1508:0] c_w_585, s_w_585;
wire [1508:0] c_w_586, s_w_586;
wire [1508:0] c_w_587, s_w_587;
wire [1508:0] c_w_588, s_w_588;
wire [1508:0] c_w_589, s_w_589;
wire [1508:0] c_w_590, s_w_590;
wire [1508:0] c_w_591, s_w_591;
wire [1508:0] c_w_592, s_w_592;
wire [1508:0] c_w_593, s_w_593;
wire [1508:0] c_w_594, s_w_594;
wire [1508:0] c_w_595, s_w_595;
wire [1508:0] c_w_596, s_w_596;
wire [1508:0] c_w_597, s_w_597;
wire [1508:0] c_w_598, s_w_598;
wire [1508:0] c_w_599, s_w_599;
wire [1508:0] c_w_600, s_w_600;
wire [1508:0] c_w_601, s_w_601;
wire [1508:0] c_w_602, s_w_602;
wire [1508:0] c_w_603, s_w_603;
wire [1508:0] c_w_604, s_w_604;
wire [1508:0] c_w_605, s_w_605;
wire [1508:0] c_w_606, s_w_606;
wire [1508:0] c_w_607, s_w_607;
wire [1508:0] c_w_608, s_w_608;
wire [1508:0] c_w_609, s_w_609;
wire [1508:0] c_w_610, s_w_610;
wire [1508:0] c_w_611, s_w_611;
wire [1508:0] c_w_612, s_w_612;
wire [1508:0] c_w_613, s_w_613;
wire [1508:0] c_w_614, s_w_614;
wire [1508:0] c_w_615, s_w_615;
wire [1508:0] c_w_616, s_w_616;
wire [1508:0] c_w_617, s_w_617;
wire [1508:0] c_w_618, s_w_618;
wire [1508:0] c_w_619, s_w_619;
wire [1508:0] c_w_620, s_w_620;
wire [1508:0] c_w_621, s_w_621;
wire [1508:0] c_w_622, s_w_622;
wire [1508:0] c_w_623, s_w_623;
wire [1508:0] c_w_624, s_w_624;
wire [1508:0] c_w_625, s_w_625;
wire [1508:0] c_w_626, s_w_626;
wire [1508:0] c_w_627, s_w_627;
wire [1508:0] c_w_628, s_w_628;
wire [1508:0] c_w_629, s_w_629;
wire [1508:0] c_w_630, s_w_630;
wire [1508:0] c_w_631, s_w_631;
wire [1508:0] c_w_632, s_w_632;
wire [1508:0] c_w_633, s_w_633;
wire [1508:0] c_w_634, s_w_634;
wire [1508:0] c_w_635, s_w_635;
wire [1508:0] c_w_636, s_w_636;
wire [1508:0] c_w_637, s_w_637;
wire [1508:0] c_w_638, s_w_638;
wire [1508:0] c_w_639, s_w_639;
wire [1508:0] c_w_640, s_w_640;
wire [1508:0] c_w_641, s_w_641;
wire [1508:0] c_w_642, s_w_642;
wire [1508:0] c_w_643, s_w_643;
wire [1508:0] c_w_644, s_w_644;
wire [1508:0] c_w_645, s_w_645;
wire [1508:0] c_w_646, s_w_646;
wire [1508:0] c_w_647, s_w_647;
wire [1508:0] c_w_648, s_w_648;
wire [1508:0] c_w_649, s_w_649;
wire [1508:0] c_w_650, s_w_650;
wire [1508:0] c_w_651, s_w_651;
wire [1508:0] c_w_652, s_w_652;
wire [1508:0] c_w_653, s_w_653;
wire [1508:0] c_w_654, s_w_654;
wire [1508:0] c_w_655, s_w_655;
wire [1508:0] c_w_656, s_w_656;
wire [1508:0] c_w_657, s_w_657;
wire [1508:0] c_w_658, s_w_658;
wire [1508:0] c_w_659, s_w_659;
wire [1508:0] c_w_660, s_w_660;
wire [1508:0] c_w_661, s_w_661;
wire [1508:0] c_w_662, s_w_662;
wire [1508:0] c_w_663, s_w_663;
wire [1508:0] c_w_664, s_w_664;
wire [1508:0] c_w_665, s_w_665;
wire [1508:0] c_w_666, s_w_666;
wire [1508:0] c_w_667, s_w_667;
wire [1508:0] c_w_668, s_w_668;
wire [1508:0] c_w_669, s_w_669;
wire [1508:0] c_w_670, s_w_670;
wire [1508:0] c_w_671, s_w_671;
wire [1508:0] c_w_672, s_w_672;
wire [1508:0] c_w_673, s_w_673;
wire [1508:0] c_w_674, s_w_674;
wire [1508:0] c_w_675, s_w_675;
wire [1508:0] c_w_676, s_w_676;
wire [1508:0] c_w_677, s_w_677;
wire [1508:0] c_w_678, s_w_678;
wire [1508:0] c_w_679, s_w_679;
wire [1508:0] c_w_680, s_w_680;
wire [1508:0] c_w_681, s_w_681;
wire [1508:0] c_w_682, s_w_682;
wire [1508:0] c_w_683, s_w_683;
wire [1508:0] c_w_684, s_w_684;
wire [1508:0] c_w_685, s_w_685;
wire [1508:0] c_w_686, s_w_686;
wire [1508:0] c_w_687, s_w_687;
wire [1508:0] c_w_688, s_w_688;
wire [1508:0] c_w_689, s_w_689;
wire [1508:0] c_w_690, s_w_690;
wire [1508:0] c_w_691, s_w_691;
wire [1508:0] c_w_692, s_w_692;
wire [1508:0] c_w_693, s_w_693;
wire [1508:0] c_w_694, s_w_694;
wire [1508:0] c_w_695, s_w_695;
wire [1508:0] c_w_696, s_w_696;
wire [1508:0] c_w_697, s_w_697;
wire [1508:0] c_w_698, s_w_698;
wire [1508:0] c_w_699, s_w_699;
wire [1508:0] c_w_700, s_w_700;
wire [1508:0] c_w_701, s_w_701;
wire [1508:0] c_w_702, s_w_702;
wire [1508:0] c_w_703, s_w_703;
wire [1508:0] c_w_704, s_w_704;
wire [1508:0] c_w_705, s_w_705;
wire [1508:0] c_w_706, s_w_706;
wire [1508:0] c_w_707, s_w_707;
wire [1508:0] c_w_708, s_w_708;
wire [1508:0] c_w_709, s_w_709;
wire [1508:0] c_w_710, s_w_710;
wire [1508:0] c_w_711, s_w_711;
wire [1508:0] c_w_712, s_w_712;
wire [1508:0] c_w_713, s_w_713;
wire [1508:0] c_w_714, s_w_714;
wire [1508:0] c_w_715, s_w_715;
wire [1508:0] c_w_716, s_w_716;
wire [1508:0] c_w_717, s_w_717;
wire [1508:0] c_w_718, s_w_718;
wire [1508:0] c_w_719, s_w_719;
wire [1508:0] c_w_720, s_w_720;
wire [1508:0] c_w_721, s_w_721;
wire [1508:0] c_w_722, s_w_722;
wire [1508:0] c_w_723, s_w_723;
wire [1508:0] c_w_724, s_w_724;
wire [1508:0] c_w_725, s_w_725;
wire [1508:0] c_w_726, s_w_726;
wire [1508:0] c_w_727, s_w_727;
wire [1508:0] c_w_728, s_w_728;
wire [1508:0] c_w_729, s_w_729;
wire [1508:0] c_w_730, s_w_730;
wire [1508:0] c_w_731, s_w_731;
wire [1508:0] c_w_732, s_w_732;
wire [1508:0] c_w_733, s_w_733;
wire [1508:0] c_w_734, s_w_734;
wire [1508:0] c_w_735, s_w_735;
wire [1508:0] c_w_736, s_w_736;
wire [1508:0] c_w_737, s_w_737;
wire [1508:0] c_w_738, s_w_738;
wire [1508:0] c_w_739, s_w_739;
wire [1508:0] c_w_740, s_w_740;
wire [1508:0] c_w_741, s_w_741;
wire [1508:0] c_w_742, s_w_742;
wire [1508:0] c_w_743, s_w_743;
wire [1508:0] c_w_744, s_w_744;
wire [1508:0] c_w_745, s_w_745;
wire [1508:0] c_w_746, s_w_746;
wire [1508:0] c_w_747, s_w_747;
wire [1508:0] c_w_748, s_w_748;
wire [1508:0] c_w_749, s_w_749;
wire [1508:0] c_w_750, s_w_750;
wire [1508:0] c_w_751, s_w_751;
wire [1508:0] c_w_752, s_w_752;
wire [1508:0] c_w_753, s_w_753;
wire [1508:0] c_w_754, s_w_754;
wire [1508:0] c_w_755, s_w_755;
wire [1508:0] c_w_756, s_w_756;
wire [1508:0] c_w_757, s_w_757;
wire [1508:0] c_w_758, s_w_758;
wire [1508:0] c_w_759, s_w_759;
wire [1508:0] c_w_760, s_w_760;
wire [1508:0] c_w_761, s_w_761;
wire [1508:0] c_w_762, s_w_762;
wire [1508:0] c_w_763, s_w_763;
wire [1508:0] c_w_764, s_w_764;
wire [1508:0] c_w_765, s_w_765;
wire [1508:0] c_w_766, s_w_766;
wire [1508:0] c_w_767, s_w_767;
wire [1508:0] c_w_768, s_w_768;
wire [1508:0] c_w_769, s_w_769;
wire [1508:0] c_w_770, s_w_770;
wire [1508:0] c_w_771, s_w_771;
wire [1508:0] c_w_772, s_w_772;
wire [1508:0] c_w_773, s_w_773;
wire [1508:0] c_w_774, s_w_774;
wire [1508:0] c_w_775, s_w_775;
wire [1508:0] c_w_776, s_w_776;
wire [1508:0] c_w_777, s_w_777;
wire [1508:0] c_w_778, s_w_778;
wire [1508:0] c_w_779, s_w_779;
wire [1508:0] c_w_780, s_w_780;
wire [1508:0] c_w_781, s_w_781;
wire [1508:0] c_w_782, s_w_782;
wire [1508:0] c_w_783, s_w_783;
wire [1508:0] c_w_784, s_w_784;
wire [1508:0] c_w_785, s_w_785;
wire [1508:0] c_w_786, s_w_786;
wire [1508:0] c_w_787, s_w_787;
wire [1508:0] c_w_788, s_w_788;
wire [1508:0] c_w_789, s_w_789;
wire [1508:0] c_w_790, s_w_790;
wire [1508:0] c_w_791, s_w_791;
wire [1508:0] c_w_792, s_w_792;
wire [1508:0] c_w_793, s_w_793;
wire [1508:0] c_w_794, s_w_794;
wire [1508:0] c_w_795, s_w_795;
wire [1508:0] c_w_796, s_w_796;
wire [1508:0] c_w_797, s_w_797;
wire [1508:0] c_w_798, s_w_798;
wire [1508:0] c_w_799, s_w_799;
wire [1508:0] c_w_800, s_w_800;
wire [1508:0] c_w_801, s_w_801;
wire [1508:0] c_w_802, s_w_802;
wire [1508:0] c_w_803, s_w_803;
wire [1508:0] c_w_804, s_w_804;
wire [1508:0] c_w_805, s_w_805;
wire [1508:0] c_w_806, s_w_806;
wire [1508:0] c_w_807, s_w_807;
wire [1508:0] c_w_808, s_w_808;
wire [1508:0] c_w_809, s_w_809;
wire [1508:0] c_w_810, s_w_810;
wire [1508:0] c_w_811, s_w_811;
wire [1508:0] c_w_812, s_w_812;
wire [1508:0] c_w_813, s_w_813;
wire [1508:0] c_w_814, s_w_814;
wire [1508:0] c_w_815, s_w_815;
wire [1508:0] c_w_816, s_w_816;
wire [1508:0] c_w_817, s_w_817;
wire [1508:0] c_w_818, s_w_818;
wire [1508:0] c_w_819, s_w_819;
wire [1508:0] c_w_820, s_w_820;
wire [1508:0] c_w_821, s_w_821;
wire [1508:0] c_w_822, s_w_822;
wire [1508:0] c_w_823, s_w_823;
wire [1508:0] c_w_824, s_w_824;
wire [1508:0] c_w_825, s_w_825;
wire [1508:0] c_w_826, s_w_826;
wire [1508:0] c_w_827, s_w_827;
wire [1508:0] c_w_828, s_w_828;
wire [1508:0] c_w_829, s_w_829;
wire [1508:0] c_w_830, s_w_830;
wire [1508:0] c_w_831, s_w_831;
wire [1508:0] c_w_832, s_w_832;
wire [1508:0] c_w_833, s_w_833;
wire [1508:0] c_w_834, s_w_834;
wire [1508:0] c_w_835, s_w_835;
wire [1508:0] c_w_836, s_w_836;
wire [1508:0] c_w_837, s_w_837;
wire [1508:0] c_w_838, s_w_838;
wire [1508:0] c_w_839, s_w_839;
wire [1508:0] c_w_840, s_w_840;
wire [1508:0] c_w_841, s_w_841;
wire [1508:0] c_w_842, s_w_842;
wire [1508:0] c_w_843, s_w_843;
wire [1508:0] c_w_844, s_w_844;
wire [1508:0] c_w_845, s_w_845;
wire [1508:0] c_w_846, s_w_846;
wire [1508:0] c_w_847, s_w_847;
wire [1508:0] c_w_848, s_w_848;
wire [1508:0] c_w_849, s_w_849;
wire [1508:0] c_w_850, s_w_850;
wire [1508:0] c_w_851, s_w_851;
wire [1508:0] c_w_852, s_w_852;
wire [1508:0] c_w_853, s_w_853;
wire [1508:0] c_w_854, s_w_854;
wire [1508:0] c_w_855, s_w_855;
wire [1508:0] c_w_856, s_w_856;
wire [1508:0] c_w_857, s_w_857;
wire [1508:0] c_w_858, s_w_858;
wire [1508:0] c_w_859, s_w_859;
wire [1508:0] c_w_860, s_w_860;
wire [1508:0] c_w_861, s_w_861;
wire [1508:0] c_w_862, s_w_862;
wire [1508:0] c_w_863, s_w_863;
wire [1508:0] c_w_864, s_w_864;
wire [1508:0] c_w_865, s_w_865;
wire [1508:0] c_w_866, s_w_866;
wire [1508:0] c_w_867, s_w_867;
wire [1508:0] c_w_868, s_w_868;
wire [1508:0] c_w_869, s_w_869;
wire [1508:0] c_w_870, s_w_870;
wire [1508:0] c_w_871, s_w_871;
wire [1508:0] c_w_872, s_w_872;
wire [1508:0] c_w_873, s_w_873;
wire [1508:0] c_w_874, s_w_874;
wire [1508:0] c_w_875, s_w_875;
wire [1508:0] c_w_876, s_w_876;
wire [1508:0] c_w_877, s_w_877;
wire [1508:0] c_w_878, s_w_878;
wire [1508:0] c_w_879, s_w_879;
wire [1508:0] c_w_880, s_w_880;
wire [1508:0] c_w_881, s_w_881;
wire [1508:0] c_w_882, s_w_882;
wire [1508:0] c_w_883, s_w_883;
wire [1508:0] c_w_884, s_w_884;
wire [1508:0] c_w_885, s_w_885;
wire [1508:0] c_w_886, s_w_886;
wire [1508:0] c_w_887, s_w_887;
wire [1508:0] c_w_888, s_w_888;
wire [1508:0] c_w_889, s_w_889;
wire [1508:0] c_w_890, s_w_890;
wire [1508:0] c_w_891, s_w_891;
wire [1508:0] c_w_892, s_w_892;
wire [1508:0] c_w_893, s_w_893;
wire [1508:0] c_w_894, s_w_894;
wire [1508:0] c_w_895, s_w_895;
wire [1508:0] c_w_896, s_w_896;
wire [1508:0] c_w_897, s_w_897;
wire [1508:0] c_w_898, s_w_898;
wire [1508:0] c_w_899, s_w_899;
wire [1508:0] c_w_900, s_w_900;
wire [1508:0] c_w_901, s_w_901;
wire [1508:0] c_w_902, s_w_902;
wire [1508:0] c_w_903, s_w_903;
wire [1508:0] c_w_904, s_w_904;
wire [1508:0] c_w_905, s_w_905;
wire [1508:0] c_w_906, s_w_906;
wire [1508:0] c_w_907, s_w_907;
wire [1508:0] c_w_908, s_w_908;
wire [1508:0] c_w_909, s_w_909;
wire [1508:0] c_w_910, s_w_910;
wire [1508:0] c_w_911, s_w_911;
wire [1508:0] c_w_912, s_w_912;
wire [1508:0] c_w_913, s_w_913;
wire [1508:0] c_w_914, s_w_914;
wire [1508:0] c_w_915, s_w_915;
wire [1508:0] c_w_916, s_w_916;
wire [1508:0] c_w_917, s_w_917;
wire [1508:0] c_w_918, s_w_918;
wire [1508:0] c_w_919, s_w_919;
wire [1508:0] c_w_920, s_w_920;
wire [1508:0] c_w_921, s_w_921;
wire [1508:0] c_w_922, s_w_922;
wire [1508:0] c_w_923, s_w_923;
wire [1508:0] c_w_924, s_w_924;
wire [1508:0] c_w_925, s_w_925;
wire [1508:0] c_w_926, s_w_926;
wire [1508:0] c_w_927, s_w_927;
wire [1508:0] c_w_928, s_w_928;
wire [1508:0] c_w_929, s_w_929;
wire [1508:0] c_w_930, s_w_930;
wire [1508:0] c_w_931, s_w_931;
wire [1508:0] c_w_932, s_w_932;
wire [1508:0] c_w_933, s_w_933;
wire [1508:0] c_w_934, s_w_934;
wire [1508:0] c_w_935, s_w_935;
wire [1508:0] c_w_936, s_w_936;
wire [1508:0] c_w_937, s_w_937;
wire [1508:0] c_w_938, s_w_938;
wire [1508:0] c_w_939, s_w_939;
wire [1508:0] c_w_940, s_w_940;
wire [1508:0] c_w_941, s_w_941;
wire [1508:0] c_w_942, s_w_942;
wire [1508:0] c_w_943, s_w_943;
wire [1508:0] c_w_944, s_w_944;
wire [1508:0] c_w_945, s_w_945;
wire [1508:0] c_w_946, s_w_946;
wire [1508:0] c_w_947, s_w_947;
wire [1508:0] c_w_948, s_w_948;
wire [1508:0] c_w_949, s_w_949;
wire [1508:0] c_w_950, s_w_950;
wire [1508:0] c_w_951, s_w_951;
wire [1508:0] c_w_952, s_w_952;
wire [1508:0] c_w_953, s_w_953;
wire [1508:0] c_w_954, s_w_954;
wire [1508:0] c_w_955, s_w_955;
wire [1508:0] c_w_956, s_w_956;
wire [1508:0] c_w_957, s_w_957;
wire [1508:0] c_w_958, s_w_958;
wire [1508:0] c_w_959, s_w_959;
wire [1508:0] c_w_960, s_w_960;
wire [1508:0] c_w_961, s_w_961;
wire [1508:0] c_w_962, s_w_962;
wire [1508:0] c_w_963, s_w_963;
wire [1508:0] c_w_964, s_w_964;
wire [1508:0] c_w_965, s_w_965;
wire [1508:0] c_w_966, s_w_966;
wire [1508:0] c_w_967, s_w_967;
wire [1508:0] c_w_968, s_w_968;
wire [1508:0] c_w_969, s_w_969;
wire [1508:0] c_w_970, s_w_970;
wire [1508:0] c_w_971, s_w_971;
wire [1508:0] c_w_972, s_w_972;
wire [1508:0] c_w_973, s_w_973;
wire [1508:0] c_w_974, s_w_974;
wire [1508:0] c_w_975, s_w_975;
wire [1508:0] c_w_976, s_w_976;
wire [1508:0] c_w_977, s_w_977;
wire [1508:0] c_w_978, s_w_978;
wire [1508:0] c_w_979, s_w_979;
wire [1508:0] c_w_980, s_w_980;
wire [1508:0] c_w_981, s_w_981;
wire [1508:0] c_w_982, s_w_982;
wire [1508:0] c_w_983, s_w_983;
wire [1508:0] c_w_984, s_w_984;
wire [1508:0] c_w_985, s_w_985;
wire [1508:0] c_w_986, s_w_986;
wire [1508:0] c_w_987, s_w_987;
wire [1508:0] c_w_988, s_w_988;
wire [1508:0] c_w_989, s_w_989;
wire [1508:0] c_w_990, s_w_990;
wire [1508:0] c_w_991, s_w_991;
wire [1508:0] c_w_992, s_w_992;
wire [1508:0] c_w_993, s_w_993;
wire [1508:0] c_w_994, s_w_994;
wire [1508:0] c_w_995, s_w_995;
wire [1508:0] c_w_996, s_w_996;
wire [1508:0] c_w_997, s_w_997;
wire [1508:0] c_w_998, s_w_998;
wire [1508:0] c_w_999, s_w_999;
wire [1508:0] c_w_1000, s_w_1000;
wire [1508:0] c_w_1001, s_w_1001;
wire [1508:0] c_w_1002, s_w_1002;
wire [1508:0] c_w_1003, s_w_1003;
wire [1508:0] c_w_1004, s_w_1004;
wire [1508:0] c_w_1005, s_w_1005;
wire [1508:0] c_w_1006, s_w_1006;
wire [1508:0] c_w_1007, s_w_1007;
wire [1508:0] c_w_1008, s_w_1008;
wire [1508:0] c_w_1009, s_w_1009;
wire [1508:0] c_w_1010, s_w_1010;
wire [1508:0] c_w_1011, s_w_1011;
wire [1508:0] c_w_1012, s_w_1012;
wire [1508:0] c_w_1013, s_w_1013;
wire [1508:0] c_w_1014, s_w_1014;
wire [1508:0] c_w_1015, s_w_1015;
wire [1508:0] c_w_1016, s_w_1016;
wire [1508:0] c_w_1017, s_w_1017;
wire [1508:0] c_w_1018, s_w_1018;
wire [1508:0] c_w_1019, s_w_1019;
wire [1508:0] c_w_1020, s_w_1020;
wire [1508:0] c_w_1021, s_w_1021;
wire [1508:0] c_w_1022, s_w_1022;
wire [1508:0] c_w_1023, s_w_1023;
wire [1508:0] c_w_1024, s_w_1024;
wire [1508:0] c_w_1025, s_w_1025;
wire [1508:0] c_w_1026, s_w_1026;
wire [1508:0] c_w_1027, s_w_1027;
wire [1508:0] c_w_1028, s_w_1028;
wire [1508:0] c_w_1029, s_w_1029;
wire [1508:0] c_w_1030, s_w_1030;
wire [1508:0] c_w_1031, s_w_1031;
wire [1508:0] c_w_1032, s_w_1032;
wire [1508:0] c_w_1033, s_w_1033;
wire [1508:0] c_w_1034, s_w_1034;
wire [1508:0] c_w_1035, s_w_1035;
wire [1508:0] c_w_1036, s_w_1036;
wire [1508:0] c_w_1037, s_w_1037;
wire [1508:0] c_w_1038, s_w_1038;
wire [1508:0] c_w_1039, s_w_1039;
wire [1508:0] c_w_1040, s_w_1040;
wire [1508:0] c_w_1041, s_w_1041;
wire [1508:0] c_w_1042, s_w_1042;
wire [1508:0] c_w_1043, s_w_1043;
wire [1508:0] c_w_1044, s_w_1044;
wire [1508:0] c_w_1045, s_w_1045;
wire [1508:0] c_w_1046, s_w_1046;
wire [1508:0] c_w_1047, s_w_1047;
wire [1508:0] c_w_1048, s_w_1048;
wire [1508:0] c_w_1049, s_w_1049;
wire [1508:0] c_w_1050, s_w_1050;
wire [1508:0] c_w_1051, s_w_1051;
wire [1508:0] c_w_1052, s_w_1052;
wire [1508:0] c_w_1053, s_w_1053;
wire [1508:0] c_w_1054, s_w_1054;
wire [1508:0] c_w_1055, s_w_1055;
wire [1508:0] c_w_1056, s_w_1056;
wire [1508:0] c_w_1057, s_w_1057;
wire [1508:0] c_w_1058, s_w_1058;
wire [1508:0] c_w_1059, s_w_1059;
wire [1508:0] c_w_1060, s_w_1060;
wire [1508:0] c_w_1061, s_w_1061;
wire [1508:0] c_w_1062, s_w_1062;
wire [1508:0] c_w_1063, s_w_1063;
wire [1508:0] c_w_1064, s_w_1064;
wire [1508:0] c_w_1065, s_w_1065;
wire [1508:0] c_w_1066, s_w_1066;
wire [1508:0] c_w_1067, s_w_1067;
wire [1508:0] c_w_1068, s_w_1068;
wire [1508:0] c_w_1069, s_w_1069;
wire [1508:0] c_w_1070, s_w_1070;
wire [1508:0] c_w_1071, s_w_1071;
wire [1508:0] c_w_1072, s_w_1072;
wire [1508:0] c_w_1073, s_w_1073;
wire [1508:0] c_w_1074, s_w_1074;
wire [1508:0] c_w_1075, s_w_1075;
wire [1508:0] c_w_1076, s_w_1076;
wire [1508:0] c_w_1077, s_w_1077;
wire [1508:0] c_w_1078, s_w_1078;
wire [1508:0] c_w_1079, s_w_1079;
wire [1508:0] c_w_1080, s_w_1080;
wire [1508:0] c_w_1081, s_w_1081;
wire [1508:0] c_w_1082, s_w_1082;
wire [1508:0] c_w_1083, s_w_1083;
wire [1508:0] c_w_1084, s_w_1084;
wire [1508:0] c_w_1085, s_w_1085;
wire [1508:0] c_w_1086, s_w_1086;
wire [1508:0] c_w_1087, s_w_1087;
wire [1508:0] c_w_1088, s_w_1088;
wire [1508:0] c_w_1089, s_w_1089;
wire [1508:0] c_w_1090, s_w_1090;
wire [1508:0] c_w_1091, s_w_1091;
wire [1508:0] c_w_1092, s_w_1092;
wire [1508:0] c_w_1093, s_w_1093;
wire [1508:0] c_w_1094, s_w_1094;
wire [1508:0] c_w_1095, s_w_1095;
wire [1508:0] c_w_1096, s_w_1096;
wire [1508:0] c_w_1097, s_w_1097;
wire [1508:0] c_w_1098, s_w_1098;
wire [1508:0] c_w_1099, s_w_1099;
wire [1508:0] c_w_1100, s_w_1100;
wire [1508:0] c_w_1101, s_w_1101;
wire [1508:0] c_w_1102, s_w_1102;
wire [1508:0] c_w_1103, s_w_1103;
wire [1508:0] c_w_1104, s_w_1104;
wire [1508:0] c_w_1105, s_w_1105;
wire [1508:0] c_w_1106, s_w_1106;
wire [1508:0] c_w_1107, s_w_1107;
wire [1508:0] c_w_1108, s_w_1108;
wire [1508:0] c_w_1109, s_w_1109;
wire [1508:0] c_w_1110, s_w_1110;
wire [1508:0] c_w_1111, s_w_1111;
wire [1508:0] c_w_1112, s_w_1112;
wire [1508:0] c_w_1113, s_w_1113;
wire [1508:0] c_w_1114, s_w_1114;
wire [1508:0] c_w_1115, s_w_1115;
wire [1508:0] c_w_1116, s_w_1116;
wire [1508:0] c_w_1117, s_w_1117;
wire [1508:0] c_w_1118, s_w_1118;
wire [1508:0] c_w_1119, s_w_1119;
wire [1508:0] c_w_1120, s_w_1120;
wire [1508:0] c_w_1121, s_w_1121;
wire [1508:0] c_w_1122, s_w_1122;
wire [1508:0] c_w_1123, s_w_1123;
wire [1508:0] c_w_1124, s_w_1124;
wire [1508:0] c_w_1125, s_w_1125;
wire [1508:0] c_w_1126, s_w_1126;
wire [1508:0] c_w_1127, s_w_1127;
wire [1508:0] c_w_1128, s_w_1128;
wire [1508:0] c_w_1129, s_w_1129;
wire [1508:0] c_w_1130, s_w_1130;
wire [1508:0] c_w_1131, s_w_1131;
wire [1508:0] c_w_1132, s_w_1132;
wire [1508:0] c_w_1133, s_w_1133;
wire [1508:0] c_w_1134, s_w_1134;
wire [1508:0] c_w_1135, s_w_1135;
wire [1508:0] c_w_1136, s_w_1136;
wire [1508:0] c_w_1137, s_w_1137;
wire [1508:0] c_w_1138, s_w_1138;
wire [1508:0] c_w_1139, s_w_1139;
wire [1508:0] c_w_1140, s_w_1140;
wire [1508:0] c_w_1141, s_w_1141;
wire [1508:0] c_w_1142, s_w_1142;
wire [1508:0] c_w_1143, s_w_1143;
wire [1508:0] c_w_1144, s_w_1144;
wire [1508:0] c_w_1145, s_w_1145;
wire [1508:0] c_w_1146, s_w_1146;
wire [1508:0] c_w_1147, s_w_1147;
wire [1508:0] c_w_1148, s_w_1148;
wire [1508:0] c_w_1149, s_w_1149;
wire [1508:0] c_w_1150, s_w_1150;
wire [1508:0] c_w_1151, s_w_1151;
wire [1508:0] c_w_1152, s_w_1152;
wire [1508:0] c_w_1153, s_w_1153;
wire [1508:0] c_w_1154, s_w_1154;
wire [1508:0] c_w_1155, s_w_1155;
wire [1508:0] c_w_1156, s_w_1156;
wire [1508:0] c_w_1157, s_w_1157;
wire [1508:0] c_w_1158, s_w_1158;
wire [1508:0] c_w_1159, s_w_1159;
wire [1508:0] c_w_1160, s_w_1160;
wire [1508:0] c_w_1161, s_w_1161;
wire [1508:0] c_w_1162, s_w_1162;
wire [1508:0] c_w_1163, s_w_1163;
wire [1508:0] c_w_1164, s_w_1164;
wire [1508:0] c_w_1165, s_w_1165;
wire [1508:0] c_w_1166, s_w_1166;
wire [1508:0] c_w_1167, s_w_1167;
wire [1508:0] c_w_1168, s_w_1168;
wire [1508:0] c_w_1169, s_w_1169;
wire [1508:0] c_w_1170, s_w_1170;
wire [1508:0] c_w_1171, s_w_1171;
wire [1508:0] c_w_1172, s_w_1172;
wire [1508:0] c_w_1173, s_w_1173;
wire [1508:0] c_w_1174, s_w_1174;
wire [1508:0] c_w_1175, s_w_1175;
wire [1508:0] c_w_1176, s_w_1176;
wire [1508:0] c_w_1177, s_w_1177;
wire [1508:0] c_w_1178, s_w_1178;
wire [1508:0] c_w_1179, s_w_1179;
wire [1508:0] c_w_1180, s_w_1180;
wire [1508:0] c_w_1181, s_w_1181;
wire [1508:0] c_w_1182, s_w_1182;
wire [1508:0] c_w_1183, s_w_1183;
wire [1508:0] c_w_1184, s_w_1184;
wire [1508:0] c_w_1185, s_w_1185;
wire [1508:0] c_w_1186, s_w_1186;
wire [1508:0] c_w_1187, s_w_1187;
wire [1508:0] c_w_1188, s_w_1188;
wire [1508:0] c_w_1189, s_w_1189;
wire [1508:0] c_w_1190, s_w_1190;
wire [1508:0] c_w_1191, s_w_1191;
wire [1508:0] c_w_1192, s_w_1192;
wire [1508:0] c_w_1193, s_w_1193;
wire [1508:0] c_w_1194, s_w_1194;
wire [1508:0] c_w_1195, s_w_1195;
wire [1508:0] c_w_1196, s_w_1196;
wire [1508:0] c_w_1197, s_w_1197;
wire [1508:0] c_w_1198, s_w_1198;
wire [1508:0] c_w_1199, s_w_1199;
wire [1508:0] c_w_1200, s_w_1200;
wire [1508:0] c_w_1201, s_w_1201;
wire [1508:0] c_w_1202, s_w_1202;
wire [1508:0] c_w_1203, s_w_1203;
wire [1508:0] c_w_1204, s_w_1204;
wire [1508:0] c_w_1205, s_w_1205;
wire [1508:0] c_w_1206, s_w_1206;
wire [1508:0] c_w_1207, s_w_1207;
wire [1508:0] c_w_1208, s_w_1208;
wire [1508:0] c_w_1209, s_w_1209;
wire [1508:0] c_w_1210, s_w_1210;
wire [1508:0] c_w_1211, s_w_1211;
wire [1508:0] c_w_1212, s_w_1212;
wire [1508:0] c_w_1213, s_w_1213;
wire [1508:0] c_w_1214, s_w_1214;
wire [1508:0] c_w_1215, s_w_1215;
wire [1508:0] c_w_1216, s_w_1216;
wire [1508:0] c_w_1217, s_w_1217;
wire [1508:0] c_w_1218, s_w_1218;
wire [1508:0] c_w_1219, s_w_1219;
wire [1508:0] c_w_1220, s_w_1220;
wire [1508:0] c_w_1221, s_w_1221;
wire [1508:0] c_w_1222, s_w_1222;
wire [1508:0] c_w_1223, s_w_1223;
wire [1508:0] c_w_1224, s_w_1224;
wire [1508:0] c_w_1225, s_w_1225;
wire [1508:0] c_w_1226, s_w_1226;
wire [1508:0] c_w_1227, s_w_1227;
wire [1508:0] c_w_1228, s_w_1228;
wire [1508:0] c_w_1229, s_w_1229;
wire [1508:0] c_w_1230, s_w_1230;
wire [1508:0] c_w_1231, s_w_1231;
wire [1508:0] c_w_1232, s_w_1232;
wire [1508:0] c_w_1233, s_w_1233;
wire [1508:0] c_w_1234, s_w_1234;
wire [1508:0] c_w_1235, s_w_1235;
wire [1508:0] c_w_1236, s_w_1236;
wire [1508:0] c_w_1237, s_w_1237;
wire [1508:0] c_w_1238, s_w_1238;
wire [1508:0] c_w_1239, s_w_1239;
wire [1508:0] c_w_1240, s_w_1240;
wire [1508:0] c_w_1241, s_w_1241;
wire [1508:0] c_w_1242, s_w_1242;
wire [1508:0] c_w_1243, s_w_1243;
wire [1508:0] c_w_1244, s_w_1244;
wire [1508:0] c_w_1245, s_w_1245;
wire [1508:0] c_w_1246, s_w_1246;
wire [1508:0] c_w_1247, s_w_1247;
wire [1508:0] c_w_1248, s_w_1248;
wire [1508:0] c_w_1249, s_w_1249;
wire [1508:0] c_w_1250, s_w_1250;
wire [1508:0] c_w_1251, s_w_1251;
wire [1508:0] c_w_1252, s_w_1252;
wire [1508:0] c_w_1253, s_w_1253;
wire [1508:0] c_w_1254, s_w_1254;
wire [1508:0] c_w_1255, s_w_1255;
wire [1508:0] c_w_1256, s_w_1256;
wire [1508:0] c_w_1257, s_w_1257;
wire [1508:0] c_w_1258, s_w_1258;
wire [1508:0] c_w_1259, s_w_1259;
wire [1508:0] c_w_1260, s_w_1260;
wire [1508:0] c_w_1261, s_w_1261;
wire [1508:0] c_w_1262, s_w_1262;
wire [1508:0] c_w_1263, s_w_1263;
wire [1508:0] c_w_1264, s_w_1264;
wire [1508:0] c_w_1265, s_w_1265;
wire [1508:0] c_w_1266, s_w_1266;
wire [1508:0] c_w_1267, s_w_1267;
wire [1508:0] c_w_1268, s_w_1268;
wire [1508:0] c_w_1269, s_w_1269;
wire [1508:0] c_w_1270, s_w_1270;
wire [1508:0] c_w_1271, s_w_1271;
wire [1508:0] c_w_1272, s_w_1272;
wire [1508:0] c_w_1273, s_w_1273;
wire [1508:0] c_w_1274, s_w_1274;
wire [1508:0] c_w_1275, s_w_1275;
wire [1508:0] c_w_1276, s_w_1276;
wire [1508:0] c_w_1277, s_w_1277;
wire [1508:0] c_w_1278, s_w_1278;
wire [1508:0] c_w_1279, s_w_1279;
wire [1508:0] c_w_1280, s_w_1280;
wire [1508:0] c_w_1281, s_w_1281;
wire [1508:0] c_w_1282, s_w_1282;
wire [1508:0] c_w_1283, s_w_1283;
wire [1508:0] c_w_1284, s_w_1284;
wire [1508:0] c_w_1285, s_w_1285;
wire [1508:0] c_w_1286, s_w_1286;
wire [1508:0] c_w_1287, s_w_1287;
wire [1508:0] c_w_1288, s_w_1288;
wire [1508:0] c_w_1289, s_w_1289;
wire [1508:0] c_w_1290, s_w_1290;
wire [1508:0] c_w_1291, s_w_1291;
wire [1508:0] c_w_1292, s_w_1292;
wire [1508:0] c_w_1293, s_w_1293;
wire [1508:0] c_w_1294, s_w_1294;
wire [1508:0] c_w_1295, s_w_1295;
wire [1508:0] c_w_1296, s_w_1296;
wire [1508:0] c_w_1297, s_w_1297;
wire [1508:0] c_w_1298, s_w_1298;
wire [1508:0] c_w_1299, s_w_1299;
wire [1508:0] c_w_1300, s_w_1300;
wire [1508:0] c_w_1301, s_w_1301;
wire [1508:0] c_w_1302, s_w_1302;
wire [1508:0] c_w_1303, s_w_1303;
wire [1508:0] c_w_1304, s_w_1304;
wire [1508:0] c_w_1305, s_w_1305;
wire [1508:0] c_w_1306, s_w_1306;
wire [1508:0] c_w_1307, s_w_1307;
wire [1508:0] c_w_1308, s_w_1308;
wire [1508:0] c_w_1309, s_w_1309;
wire [1508:0] c_w_1310, s_w_1310;
wire [1508:0] c_w_1311, s_w_1311;
wire [1508:0] c_w_1312, s_w_1312;
wire [1508:0] c_w_1313, s_w_1313;
wire [1508:0] c_w_1314, s_w_1314;
wire [1508:0] c_w_1315, s_w_1315;
wire [1508:0] c_w_1316, s_w_1316;
wire [1508:0] c_w_1317, s_w_1317;
wire [1508:0] c_w_1318, s_w_1318;
wire [1508:0] c_w_1319, s_w_1319;
wire [1508:0] c_w_1320, s_w_1320;
wire [1508:0] c_w_1321, s_w_1321;
wire [1508:0] c_w_1322, s_w_1322;
wire [1508:0] c_w_1323, s_w_1323;
wire [1508:0] c_w_1324, s_w_1324;
wire [1508:0] c_w_1325, s_w_1325;
wire [1508:0] c_w_1326, s_w_1326;
wire [1508:0] c_w_1327, s_w_1327;
wire [1508:0] c_w_1328, s_w_1328;
wire [1508:0] c_w_1329, s_w_1329;
wire [1508:0] c_w_1330, s_w_1330;
wire [1508:0] c_w_1331, s_w_1331;
wire [1508:0] c_w_1332, s_w_1332;
wire [1508:0] c_w_1333, s_w_1333;
wire [1508:0] c_w_1334, s_w_1334;
wire [1508:0] c_w_1335, s_w_1335;
wire [1508:0] c_w_1336, s_w_1336;
wire [1508:0] c_w_1337, s_w_1337;
wire [1508:0] c_w_1338, s_w_1338;
wire [1508:0] c_w_1339, s_w_1339;
wire [1508:0] c_w_1340, s_w_1340;
wire [1508:0] c_w_1341, s_w_1341;
wire [1508:0] c_w_1342, s_w_1342;
wire [1508:0] c_w_1343, s_w_1343;
wire [1508:0] c_w_1344, s_w_1344;
wire [1508:0] c_w_1345, s_w_1345;
wire [1508:0] c_w_1346, s_w_1346;
wire [1508:0] c_w_1347, s_w_1347;
wire [1508:0] c_w_1348, s_w_1348;
wire [1508:0] c_w_1349, s_w_1349;
wire [1508:0] c_w_1350, s_w_1350;
wire [1508:0] c_w_1351, s_w_1351;
wire [1508:0] c_w_1352, s_w_1352;
wire [1508:0] c_w_1353, s_w_1353;
wire [1508:0] c_w_1354, s_w_1354;
wire [1508:0] c_w_1355, s_w_1355;
wire [1508:0] c_w_1356, s_w_1356;
wire [1508:0] c_w_1357, s_w_1357;
wire [1508:0] c_w_1358, s_w_1358;
wire [1508:0] c_w_1359, s_w_1359;
wire [1508:0] c_w_1360, s_w_1360;
wire [1508:0] c_w_1361, s_w_1361;
wire [1508:0] c_w_1362, s_w_1362;
wire [1508:0] c_w_1363, s_w_1363;
wire [1508:0] c_w_1364, s_w_1364;
wire [1508:0] c_w_1365, s_w_1365;
wire [1508:0] c_w_1366, s_w_1366;
wire [1508:0] c_w_1367, s_w_1367;
wire [1508:0] c_w_1368, s_w_1368;
wire [1508:0] c_w_1369, s_w_1369;
wire [1508:0] c_w_1370, s_w_1370;
wire [1508:0] c_w_1371, s_w_1371;
wire [1508:0] c_w_1372, s_w_1372;
wire [1508:0] c_w_1373, s_w_1373;
wire [1508:0] c_w_1374, s_w_1374;
wire [1508:0] c_w_1375, s_w_1375;
wire [1508:0] c_w_1376, s_w_1376;
wire [1508:0] c_w_1377, s_w_1377;
wire [1508:0] c_w_1378, s_w_1378;
wire [1508:0] c_w_1379, s_w_1379;
wire [1508:0] c_w_1380, s_w_1380;
wire [1508:0] c_w_1381, s_w_1381;
wire [1508:0] c_w_1382, s_w_1382;
wire [1508:0] c_w_1383, s_w_1383;
wire [1508:0] c_w_1384, s_w_1384;
wire [1508:0] c_w_1385, s_w_1385;
wire [1508:0] c_w_1386, s_w_1386;
wire [1508:0] c_w_1387, s_w_1387;
wire [1508:0] c_w_1388, s_w_1388;
wire [1508:0] c_w_1389, s_w_1389;
wire [1508:0] c_w_1390, s_w_1390;
wire [1508:0] c_w_1391, s_w_1391;
wire [1508:0] c_w_1392, s_w_1392;
wire [1508:0] c_w_1393, s_w_1393;
wire [1508:0] c_w_1394, s_w_1394;
wire [1508:0] c_w_1395, s_w_1395;
wire [1508:0] c_w_1396, s_w_1396;
wire [1508:0] c_w_1397, s_w_1397;
wire [1508:0] c_w_1398, s_w_1398;
wire [1508:0] c_w_1399, s_w_1399;
wire [1508:0] c_w_1400, s_w_1400;
wire [1508:0] c_w_1401, s_w_1401;
wire [1508:0] c_w_1402, s_w_1402;
wire [1508:0] c_w_1403, s_w_1403;
wire [1508:0] c_w_1404, s_w_1404;
wire [1508:0] c_w_1405, s_w_1405;
wire [1508:0] c_w_1406, s_w_1406;
wire [1508:0] c_w_1407, s_w_1407;
wire [1508:0] c_w_1408, s_w_1408;
wire [1508:0] c_w_1409, s_w_1409;
wire [1508:0] c_w_1410, s_w_1410;
wire [1508:0] c_w_1411, s_w_1411;
wire [1508:0] c_w_1412, s_w_1412;
wire [1508:0] c_w_1413, s_w_1413;
wire [1508:0] c_w_1414, s_w_1414;
wire [1508:0] c_w_1415, s_w_1415;
wire [1508:0] c_w_1416, s_w_1416;
wire [1508:0] c_w_1417, s_w_1417;
wire [1508:0] c_w_1418, s_w_1418;
wire [1508:0] c_w_1419, s_w_1419;
wire [1508:0] c_w_1420, s_w_1420;
wire [1508:0] c_w_1421, s_w_1421;
wire [1508:0] c_w_1422, s_w_1422;
wire [1508:0] c_w_1423, s_w_1423;
wire [1508:0] c_w_1424, s_w_1424;
wire [1508:0] c_w_1425, s_w_1425;
wire [1508:0] c_w_1426, s_w_1426;
wire [1508:0] c_w_1427, s_w_1427;
wire [1508:0] c_w_1428, s_w_1428;
wire [1508:0] c_w_1429, s_w_1429;
wire [1508:0] c_w_1430, s_w_1430;
wire [1508:0] c_w_1431, s_w_1431;
wire [1508:0] c_w_1432, s_w_1432;
wire [1508:0] c_w_1433, s_w_1433;
wire [1508:0] c_w_1434, s_w_1434;
wire [1508:0] c_w_1435, s_w_1435;
wire [1508:0] c_w_1436, s_w_1436;
wire [1508:0] c_w_1437, s_w_1437;
wire [1508:0] c_w_1438, s_w_1438;
wire [1508:0] c_w_1439, s_w_1439;
wire [1508:0] c_w_1440, s_w_1440;
wire [1508:0] c_w_1441, s_w_1441;
wire [1508:0] c_w_1442, s_w_1442;
wire [1508:0] c_w_1443, s_w_1443;
wire [1508:0] c_w_1444, s_w_1444;
wire [1508:0] c_w_1445, s_w_1445;
wire [1508:0] c_w_1446, s_w_1446;
wire [1508:0] c_w_1447, s_w_1447;
wire [1508:0] c_w_1448, s_w_1448;
wire [1508:0] c_w_1449, s_w_1449;
wire [1508:0] c_w_1450, s_w_1450;
wire [1508:0] c_w_1451, s_w_1451;
wire [1508:0] c_w_1452, s_w_1452;
wire [1508:0] c_w_1453, s_w_1453;
wire [1508:0] c_w_1454, s_w_1454;
wire [1508:0] c_w_1455, s_w_1455;
wire [1508:0] c_w_1456, s_w_1456;
wire [1508:0] c_w_1457, s_w_1457;
wire [1508:0] c_w_1458, s_w_1458;
wire [1508:0] c_w_1459, s_w_1459;
wire [1508:0] c_w_1460, s_w_1460;
wire [1508:0] c_w_1461, s_w_1461;
wire [1508:0] c_w_1462, s_w_1462;
wire [1508:0] c_w_1463, s_w_1463;
wire [1508:0] c_w_1464, s_w_1464;
wire [1508:0] c_w_1465, s_w_1465;
wire [1508:0] c_w_1466, s_w_1466;
wire [1508:0] c_w_1467, s_w_1467;
wire [1508:0] c_w_1468, s_w_1468;
wire [1508:0] c_w_1469, s_w_1469;
wire [1508:0] c_w_1470, s_w_1470;
wire [1508:0] c_w_1471, s_w_1471;
wire [1508:0] c_w_1472, s_w_1472;
wire [1508:0] c_w_1473, s_w_1473;
wire [1508:0] c_w_1474, s_w_1474;
wire [1508:0] c_w_1475, s_w_1475;
wire [1508:0] c_w_1476, s_w_1476;
wire [1508:0] c_w_1477, s_w_1477;
wire [1508:0] c_w_1478, s_w_1478;
wire [1508:0] c_w_1479, s_w_1479;
wire [1508:0] c_w_1480, s_w_1480;
wire [1508:0] c_w_1481, s_w_1481;
wire [1508:0] c_w_1482, s_w_1482;
wire [1508:0] c_w_1483, s_w_1483;
wire [1508:0] c_w_1484, s_w_1484;
wire [1508:0] c_w_1485, s_w_1485;
wire [1508:0] c_w_1486, s_w_1486;
wire [1508:0] c_w_1487, s_w_1487;
wire [1508:0] c_w_1488, s_w_1488;
wire [1508:0] c_w_1489, s_w_1489;
wire [1508:0] c_w_1490, s_w_1490;
wire [1508:0] c_w_1491, s_w_1491;
wire [1508:0] c_w_1492, s_w_1492;
wire [1508:0] c_w_1493, s_w_1493;
wire [1508:0] c_w_1494, s_w_1494;
wire [1508:0] c_w_1495, s_w_1495;
wire [1508:0] c_w_1496, s_w_1496;
wire [1508:0] c_w_1497, s_w_1497;
wire [1508:0] c_w_1498, s_w_1498;
wire [1508:0] c_w_1499, s_w_1499;
wire [1508:0] c_w_1500, s_w_1500;
wire [1508:0] c_w_1501, s_w_1501;
wire [1508:0] c_w_1502, s_w_1502;
wire [1508:0] c_w_1503, s_w_1503;
wire [1508:0] c_w_1504, s_w_1504;
wire [1508:0] c_w_1505, s_w_1505;
wire [1508:0] c_w_1506, s_w_1506;
wire [1508:0] c_w_1507, s_w_1507;
wire [1508:0] c_w_1508, s_w_1508;
    
AND_array_1509 AND_array_1509_c0({a_c[1508:0]},p_prime[0],c_w_0);
AND_array_1509 AND_array_1509_s0({a_s[1508:0]},p_prime[0],s_w_0);
AND_array_1509 AND_array_1509_c1({a_c[1507:0],1'd0},p_prime[1],c_w_1);
AND_array_1509 AND_array_1509_s1({a_s[1507:0],1'd0},p_prime[1],s_w_1);
AND_array_1509 AND_array_1509_c2({a_c[1506:0],2'd0},p_prime[2],c_w_2);
AND_array_1509 AND_array_1509_s2({a_s[1506:0],2'd0},p_prime[2],s_w_2);
AND_array_1509 AND_array_1509_c3({a_c[1505:0],3'd0},p_prime[3],c_w_3);
AND_array_1509 AND_array_1509_s3({a_s[1505:0],3'd0},p_prime[3],s_w_3);
AND_array_1509 AND_array_1509_c4({a_c[1504:0],4'd0},p_prime[4],c_w_4);
AND_array_1509 AND_array_1509_s4({a_s[1504:0],4'd0},p_prime[4],s_w_4);
AND_array_1509 AND_array_1509_c5({a_c[1503:0],5'd0},p_prime[5],c_w_5);
AND_array_1509 AND_array_1509_s5({a_s[1503:0],5'd0},p_prime[5],s_w_5);
AND_array_1509 AND_array_1509_c6({a_c[1502:0],6'd0},p_prime[6],c_w_6);
AND_array_1509 AND_array_1509_s6({a_s[1502:0],6'd0},p_prime[6],s_w_6);
AND_array_1509 AND_array_1509_c7({a_c[1501:0],7'd0},p_prime[7],c_w_7);
AND_array_1509 AND_array_1509_s7({a_s[1501:0],7'd0},p_prime[7],s_w_7);
AND_array_1509 AND_array_1509_c8({a_c[1500:0],8'd0},p_prime[8],c_w_8);
AND_array_1509 AND_array_1509_s8({a_s[1500:0],8'd0},p_prime[8],s_w_8);
AND_array_1509 AND_array_1509_c9({a_c[1499:0],9'd0},p_prime[9],c_w_9);
AND_array_1509 AND_array_1509_s9({a_s[1499:0],9'd0},p_prime[9],s_w_9);
AND_array_1509 AND_array_1509_c10({a_c[1498:0],10'd0},p_prime[10],c_w_10);
AND_array_1509 AND_array_1509_s10({a_s[1498:0],10'd0},p_prime[10],s_w_10);
AND_array_1509 AND_array_1509_c11({a_c[1497:0],11'd0},p_prime[11],c_w_11);
AND_array_1509 AND_array_1509_s11({a_s[1497:0],11'd0},p_prime[11],s_w_11);
AND_array_1509 AND_array_1509_c12({a_c[1496:0],12'd0},p_prime[12],c_w_12);
AND_array_1509 AND_array_1509_s12({a_s[1496:0],12'd0},p_prime[12],s_w_12);
AND_array_1509 AND_array_1509_c13({a_c[1495:0],13'd0},p_prime[13],c_w_13);
AND_array_1509 AND_array_1509_s13({a_s[1495:0],13'd0},p_prime[13],s_w_13);
AND_array_1509 AND_array_1509_c14({a_c[1494:0],14'd0},p_prime[14],c_w_14);
AND_array_1509 AND_array_1509_s14({a_s[1494:0],14'd0},p_prime[14],s_w_14);
AND_array_1509 AND_array_1509_c15({a_c[1493:0],15'd0},p_prime[15],c_w_15);
AND_array_1509 AND_array_1509_s15({a_s[1493:0],15'd0},p_prime[15],s_w_15);
AND_array_1509 AND_array_1509_c16({a_c[1492:0],16'd0},p_prime[16],c_w_16);
AND_array_1509 AND_array_1509_s16({a_s[1492:0],16'd0},p_prime[16],s_w_16);
AND_array_1509 AND_array_1509_c17({a_c[1491:0],17'd0},p_prime[17],c_w_17);
AND_array_1509 AND_array_1509_s17({a_s[1491:0],17'd0},p_prime[17],s_w_17);
AND_array_1509 AND_array_1509_c18({a_c[1490:0],18'd0},p_prime[18],c_w_18);
AND_array_1509 AND_array_1509_s18({a_s[1490:0],18'd0},p_prime[18],s_w_18);
AND_array_1509 AND_array_1509_c19({a_c[1489:0],19'd0},p_prime[19],c_w_19);
AND_array_1509 AND_array_1509_s19({a_s[1489:0],19'd0},p_prime[19],s_w_19);
AND_array_1509 AND_array_1509_c20({a_c[1488:0],20'd0},p_prime[20],c_w_20);
AND_array_1509 AND_array_1509_s20({a_s[1488:0],20'd0},p_prime[20],s_w_20);
AND_array_1509 AND_array_1509_c21({a_c[1487:0],21'd0},p_prime[21],c_w_21);
AND_array_1509 AND_array_1509_s21({a_s[1487:0],21'd0},p_prime[21],s_w_21);
AND_array_1509 AND_array_1509_c22({a_c[1486:0],22'd0},p_prime[22],c_w_22);
AND_array_1509 AND_array_1509_s22({a_s[1486:0],22'd0},p_prime[22],s_w_22);
AND_array_1509 AND_array_1509_c23({a_c[1485:0],23'd0},p_prime[23],c_w_23);
AND_array_1509 AND_array_1509_s23({a_s[1485:0],23'd0},p_prime[23],s_w_23);
AND_array_1509 AND_array_1509_c24({a_c[1484:0],24'd0},p_prime[24],c_w_24);
AND_array_1509 AND_array_1509_s24({a_s[1484:0],24'd0},p_prime[24],s_w_24);
AND_array_1509 AND_array_1509_c25({a_c[1483:0],25'd0},p_prime[25],c_w_25);
AND_array_1509 AND_array_1509_s25({a_s[1483:0],25'd0},p_prime[25],s_w_25);
AND_array_1509 AND_array_1509_c26({a_c[1482:0],26'd0},p_prime[26],c_w_26);
AND_array_1509 AND_array_1509_s26({a_s[1482:0],26'd0},p_prime[26],s_w_26);
AND_array_1509 AND_array_1509_c27({a_c[1481:0],27'd0},p_prime[27],c_w_27);
AND_array_1509 AND_array_1509_s27({a_s[1481:0],27'd0},p_prime[27],s_w_27);
AND_array_1509 AND_array_1509_c28({a_c[1480:0],28'd0},p_prime[28],c_w_28);
AND_array_1509 AND_array_1509_s28({a_s[1480:0],28'd0},p_prime[28],s_w_28);
AND_array_1509 AND_array_1509_c29({a_c[1479:0],29'd0},p_prime[29],c_w_29);
AND_array_1509 AND_array_1509_s29({a_s[1479:0],29'd0},p_prime[29],s_w_29);
AND_array_1509 AND_array_1509_c30({a_c[1478:0],30'd0},p_prime[30],c_w_30);
AND_array_1509 AND_array_1509_s30({a_s[1478:0],30'd0},p_prime[30],s_w_30);
AND_array_1509 AND_array_1509_c31({a_c[1477:0],31'd0},p_prime[31],c_w_31);
AND_array_1509 AND_array_1509_s31({a_s[1477:0],31'd0},p_prime[31],s_w_31);
AND_array_1509 AND_array_1509_c32({a_c[1476:0],32'd0},p_prime[32],c_w_32);
AND_array_1509 AND_array_1509_s32({a_s[1476:0],32'd0},p_prime[32],s_w_32);
AND_array_1509 AND_array_1509_c33({a_c[1475:0],33'd0},p_prime[33],c_w_33);
AND_array_1509 AND_array_1509_s33({a_s[1475:0],33'd0},p_prime[33],s_w_33);
AND_array_1509 AND_array_1509_c34({a_c[1474:0],34'd0},p_prime[34],c_w_34);
AND_array_1509 AND_array_1509_s34({a_s[1474:0],34'd0},p_prime[34],s_w_34);
AND_array_1509 AND_array_1509_c35({a_c[1473:0],35'd0},p_prime[35],c_w_35);
AND_array_1509 AND_array_1509_s35({a_s[1473:0],35'd0},p_prime[35],s_w_35);
AND_array_1509 AND_array_1509_c36({a_c[1472:0],36'd0},p_prime[36],c_w_36);
AND_array_1509 AND_array_1509_s36({a_s[1472:0],36'd0},p_prime[36],s_w_36);
AND_array_1509 AND_array_1509_c37({a_c[1471:0],37'd0},p_prime[37],c_w_37);
AND_array_1509 AND_array_1509_s37({a_s[1471:0],37'd0},p_prime[37],s_w_37);
AND_array_1509 AND_array_1509_c38({a_c[1470:0],38'd0},p_prime[38],c_w_38);
AND_array_1509 AND_array_1509_s38({a_s[1470:0],38'd0},p_prime[38],s_w_38);
AND_array_1509 AND_array_1509_c39({a_c[1469:0],39'd0},p_prime[39],c_w_39);
AND_array_1509 AND_array_1509_s39({a_s[1469:0],39'd0},p_prime[39],s_w_39);
AND_array_1509 AND_array_1509_c40({a_c[1468:0],40'd0},p_prime[40],c_w_40);
AND_array_1509 AND_array_1509_s40({a_s[1468:0],40'd0},p_prime[40],s_w_40);
AND_array_1509 AND_array_1509_c41({a_c[1467:0],41'd0},p_prime[41],c_w_41);
AND_array_1509 AND_array_1509_s41({a_s[1467:0],41'd0},p_prime[41],s_w_41);
AND_array_1509 AND_array_1509_c42({a_c[1466:0],42'd0},p_prime[42],c_w_42);
AND_array_1509 AND_array_1509_s42({a_s[1466:0],42'd0},p_prime[42],s_w_42);
AND_array_1509 AND_array_1509_c43({a_c[1465:0],43'd0},p_prime[43],c_w_43);
AND_array_1509 AND_array_1509_s43({a_s[1465:0],43'd0},p_prime[43],s_w_43);
AND_array_1509 AND_array_1509_c44({a_c[1464:0],44'd0},p_prime[44],c_w_44);
AND_array_1509 AND_array_1509_s44({a_s[1464:0],44'd0},p_prime[44],s_w_44);
AND_array_1509 AND_array_1509_c45({a_c[1463:0],45'd0},p_prime[45],c_w_45);
AND_array_1509 AND_array_1509_s45({a_s[1463:0],45'd0},p_prime[45],s_w_45);
AND_array_1509 AND_array_1509_c46({a_c[1462:0],46'd0},p_prime[46],c_w_46);
AND_array_1509 AND_array_1509_s46({a_s[1462:0],46'd0},p_prime[46],s_w_46);
AND_array_1509 AND_array_1509_c47({a_c[1461:0],47'd0},p_prime[47],c_w_47);
AND_array_1509 AND_array_1509_s47({a_s[1461:0],47'd0},p_prime[47],s_w_47);
AND_array_1509 AND_array_1509_c48({a_c[1460:0],48'd0},p_prime[48],c_w_48);
AND_array_1509 AND_array_1509_s48({a_s[1460:0],48'd0},p_prime[48],s_w_48);
AND_array_1509 AND_array_1509_c49({a_c[1459:0],49'd0},p_prime[49],c_w_49);
AND_array_1509 AND_array_1509_s49({a_s[1459:0],49'd0},p_prime[49],s_w_49);
AND_array_1509 AND_array_1509_c50({a_c[1458:0],50'd0},p_prime[50],c_w_50);
AND_array_1509 AND_array_1509_s50({a_s[1458:0],50'd0},p_prime[50],s_w_50);
AND_array_1509 AND_array_1509_c51({a_c[1457:0],51'd0},p_prime[51],c_w_51);
AND_array_1509 AND_array_1509_s51({a_s[1457:0],51'd0},p_prime[51],s_w_51);
AND_array_1509 AND_array_1509_c52({a_c[1456:0],52'd0},p_prime[52],c_w_52);
AND_array_1509 AND_array_1509_s52({a_s[1456:0],52'd0},p_prime[52],s_w_52);
AND_array_1509 AND_array_1509_c53({a_c[1455:0],53'd0},p_prime[53],c_w_53);
AND_array_1509 AND_array_1509_s53({a_s[1455:0],53'd0},p_prime[53],s_w_53);
AND_array_1509 AND_array_1509_c54({a_c[1454:0],54'd0},p_prime[54],c_w_54);
AND_array_1509 AND_array_1509_s54({a_s[1454:0],54'd0},p_prime[54],s_w_54);
AND_array_1509 AND_array_1509_c55({a_c[1453:0],55'd0},p_prime[55],c_w_55);
AND_array_1509 AND_array_1509_s55({a_s[1453:0],55'd0},p_prime[55],s_w_55);
AND_array_1509 AND_array_1509_c56({a_c[1452:0],56'd0},p_prime[56],c_w_56);
AND_array_1509 AND_array_1509_s56({a_s[1452:0],56'd0},p_prime[56],s_w_56);
AND_array_1509 AND_array_1509_c57({a_c[1451:0],57'd0},p_prime[57],c_w_57);
AND_array_1509 AND_array_1509_s57({a_s[1451:0],57'd0},p_prime[57],s_w_57);
AND_array_1509 AND_array_1509_c58({a_c[1450:0],58'd0},p_prime[58],c_w_58);
AND_array_1509 AND_array_1509_s58({a_s[1450:0],58'd0},p_prime[58],s_w_58);
AND_array_1509 AND_array_1509_c59({a_c[1449:0],59'd0},p_prime[59],c_w_59);
AND_array_1509 AND_array_1509_s59({a_s[1449:0],59'd0},p_prime[59],s_w_59);
AND_array_1509 AND_array_1509_c60({a_c[1448:0],60'd0},p_prime[60],c_w_60);
AND_array_1509 AND_array_1509_s60({a_s[1448:0],60'd0},p_prime[60],s_w_60);
AND_array_1509 AND_array_1509_c61({a_c[1447:0],61'd0},p_prime[61],c_w_61);
AND_array_1509 AND_array_1509_s61({a_s[1447:0],61'd0},p_prime[61],s_w_61);
AND_array_1509 AND_array_1509_c62({a_c[1446:0],62'd0},p_prime[62],c_w_62);
AND_array_1509 AND_array_1509_s62({a_s[1446:0],62'd0},p_prime[62],s_w_62);
AND_array_1509 AND_array_1509_c63({a_c[1445:0],63'd0},p_prime[63],c_w_63);
AND_array_1509 AND_array_1509_s63({a_s[1445:0],63'd0},p_prime[63],s_w_63);
AND_array_1509 AND_array_1509_c64({a_c[1444:0],64'd0},p_prime[64],c_w_64);
AND_array_1509 AND_array_1509_s64({a_s[1444:0],64'd0},p_prime[64],s_w_64);
AND_array_1509 AND_array_1509_c65({a_c[1443:0],65'd0},p_prime[65],c_w_65);
AND_array_1509 AND_array_1509_s65({a_s[1443:0],65'd0},p_prime[65],s_w_65);
AND_array_1509 AND_array_1509_c66({a_c[1442:0],66'd0},p_prime[66],c_w_66);
AND_array_1509 AND_array_1509_s66({a_s[1442:0],66'd0},p_prime[66],s_w_66);
AND_array_1509 AND_array_1509_c67({a_c[1441:0],67'd0},p_prime[67],c_w_67);
AND_array_1509 AND_array_1509_s67({a_s[1441:0],67'd0},p_prime[67],s_w_67);
AND_array_1509 AND_array_1509_c68({a_c[1440:0],68'd0},p_prime[68],c_w_68);
AND_array_1509 AND_array_1509_s68({a_s[1440:0],68'd0},p_prime[68],s_w_68);
AND_array_1509 AND_array_1509_c69({a_c[1439:0],69'd0},p_prime[69],c_w_69);
AND_array_1509 AND_array_1509_s69({a_s[1439:0],69'd0},p_prime[69],s_w_69);
AND_array_1509 AND_array_1509_c70({a_c[1438:0],70'd0},p_prime[70],c_w_70);
AND_array_1509 AND_array_1509_s70({a_s[1438:0],70'd0},p_prime[70],s_w_70);
AND_array_1509 AND_array_1509_c71({a_c[1437:0],71'd0},p_prime[71],c_w_71);
AND_array_1509 AND_array_1509_s71({a_s[1437:0],71'd0},p_prime[71],s_w_71);
AND_array_1509 AND_array_1509_c72({a_c[1436:0],72'd0},p_prime[72],c_w_72);
AND_array_1509 AND_array_1509_s72({a_s[1436:0],72'd0},p_prime[72],s_w_72);
AND_array_1509 AND_array_1509_c73({a_c[1435:0],73'd0},p_prime[73],c_w_73);
AND_array_1509 AND_array_1509_s73({a_s[1435:0],73'd0},p_prime[73],s_w_73);
AND_array_1509 AND_array_1509_c74({a_c[1434:0],74'd0},p_prime[74],c_w_74);
AND_array_1509 AND_array_1509_s74({a_s[1434:0],74'd0},p_prime[74],s_w_74);
AND_array_1509 AND_array_1509_c75({a_c[1433:0],75'd0},p_prime[75],c_w_75);
AND_array_1509 AND_array_1509_s75({a_s[1433:0],75'd0},p_prime[75],s_w_75);
AND_array_1509 AND_array_1509_c76({a_c[1432:0],76'd0},p_prime[76],c_w_76);
AND_array_1509 AND_array_1509_s76({a_s[1432:0],76'd0},p_prime[76],s_w_76);
AND_array_1509 AND_array_1509_c77({a_c[1431:0],77'd0},p_prime[77],c_w_77);
AND_array_1509 AND_array_1509_s77({a_s[1431:0],77'd0},p_prime[77],s_w_77);
AND_array_1509 AND_array_1509_c78({a_c[1430:0],78'd0},p_prime[78],c_w_78);
AND_array_1509 AND_array_1509_s78({a_s[1430:0],78'd0},p_prime[78],s_w_78);
AND_array_1509 AND_array_1509_c79({a_c[1429:0],79'd0},p_prime[79],c_w_79);
AND_array_1509 AND_array_1509_s79({a_s[1429:0],79'd0},p_prime[79],s_w_79);
AND_array_1509 AND_array_1509_c80({a_c[1428:0],80'd0},p_prime[80],c_w_80);
AND_array_1509 AND_array_1509_s80({a_s[1428:0],80'd0},p_prime[80],s_w_80);
AND_array_1509 AND_array_1509_c81({a_c[1427:0],81'd0},p_prime[81],c_w_81);
AND_array_1509 AND_array_1509_s81({a_s[1427:0],81'd0},p_prime[81],s_w_81);
AND_array_1509 AND_array_1509_c82({a_c[1426:0],82'd0},p_prime[82],c_w_82);
AND_array_1509 AND_array_1509_s82({a_s[1426:0],82'd0},p_prime[82],s_w_82);
AND_array_1509 AND_array_1509_c83({a_c[1425:0],83'd0},p_prime[83],c_w_83);
AND_array_1509 AND_array_1509_s83({a_s[1425:0],83'd0},p_prime[83],s_w_83);
AND_array_1509 AND_array_1509_c84({a_c[1424:0],84'd0},p_prime[84],c_w_84);
AND_array_1509 AND_array_1509_s84({a_s[1424:0],84'd0},p_prime[84],s_w_84);
AND_array_1509 AND_array_1509_c85({a_c[1423:0],85'd0},p_prime[85],c_w_85);
AND_array_1509 AND_array_1509_s85({a_s[1423:0],85'd0},p_prime[85],s_w_85);
AND_array_1509 AND_array_1509_c86({a_c[1422:0],86'd0},p_prime[86],c_w_86);
AND_array_1509 AND_array_1509_s86({a_s[1422:0],86'd0},p_prime[86],s_w_86);
AND_array_1509 AND_array_1509_c87({a_c[1421:0],87'd0},p_prime[87],c_w_87);
AND_array_1509 AND_array_1509_s87({a_s[1421:0],87'd0},p_prime[87],s_w_87);
AND_array_1509 AND_array_1509_c88({a_c[1420:0],88'd0},p_prime[88],c_w_88);
AND_array_1509 AND_array_1509_s88({a_s[1420:0],88'd0},p_prime[88],s_w_88);
AND_array_1509 AND_array_1509_c89({a_c[1419:0],89'd0},p_prime[89],c_w_89);
AND_array_1509 AND_array_1509_s89({a_s[1419:0],89'd0},p_prime[89],s_w_89);
AND_array_1509 AND_array_1509_c90({a_c[1418:0],90'd0},p_prime[90],c_w_90);
AND_array_1509 AND_array_1509_s90({a_s[1418:0],90'd0},p_prime[90],s_w_90);
AND_array_1509 AND_array_1509_c91({a_c[1417:0],91'd0},p_prime[91],c_w_91);
AND_array_1509 AND_array_1509_s91({a_s[1417:0],91'd0},p_prime[91],s_w_91);
AND_array_1509 AND_array_1509_c92({a_c[1416:0],92'd0},p_prime[92],c_w_92);
AND_array_1509 AND_array_1509_s92({a_s[1416:0],92'd0},p_prime[92],s_w_92);
AND_array_1509 AND_array_1509_c93({a_c[1415:0],93'd0},p_prime[93],c_w_93);
AND_array_1509 AND_array_1509_s93({a_s[1415:0],93'd0},p_prime[93],s_w_93);
AND_array_1509 AND_array_1509_c94({a_c[1414:0],94'd0},p_prime[94],c_w_94);
AND_array_1509 AND_array_1509_s94({a_s[1414:0],94'd0},p_prime[94],s_w_94);
AND_array_1509 AND_array_1509_c95({a_c[1413:0],95'd0},p_prime[95],c_w_95);
AND_array_1509 AND_array_1509_s95({a_s[1413:0],95'd0},p_prime[95],s_w_95);
AND_array_1509 AND_array_1509_c96({a_c[1412:0],96'd0},p_prime[96],c_w_96);
AND_array_1509 AND_array_1509_s96({a_s[1412:0],96'd0},p_prime[96],s_w_96);
AND_array_1509 AND_array_1509_c97({a_c[1411:0],97'd0},p_prime[97],c_w_97);
AND_array_1509 AND_array_1509_s97({a_s[1411:0],97'd0},p_prime[97],s_w_97);
AND_array_1509 AND_array_1509_c98({a_c[1410:0],98'd0},p_prime[98],c_w_98);
AND_array_1509 AND_array_1509_s98({a_s[1410:0],98'd0},p_prime[98],s_w_98);
AND_array_1509 AND_array_1509_c99({a_c[1409:0],99'd0},p_prime[99],c_w_99);
AND_array_1509 AND_array_1509_s99({a_s[1409:0],99'd0},p_prime[99],s_w_99);
AND_array_1509 AND_array_1509_c100({a_c[1408:0],100'd0},p_prime[100],c_w_100);
AND_array_1509 AND_array_1509_s100({a_s[1408:0],100'd0},p_prime[100],s_w_100);
AND_array_1509 AND_array_1509_c101({a_c[1407:0],101'd0},p_prime[101],c_w_101);
AND_array_1509 AND_array_1509_s101({a_s[1407:0],101'd0},p_prime[101],s_w_101);
AND_array_1509 AND_array_1509_c102({a_c[1406:0],102'd0},p_prime[102],c_w_102);
AND_array_1509 AND_array_1509_s102({a_s[1406:0],102'd0},p_prime[102],s_w_102);
AND_array_1509 AND_array_1509_c103({a_c[1405:0],103'd0},p_prime[103],c_w_103);
AND_array_1509 AND_array_1509_s103({a_s[1405:0],103'd0},p_prime[103],s_w_103);
AND_array_1509 AND_array_1509_c104({a_c[1404:0],104'd0},p_prime[104],c_w_104);
AND_array_1509 AND_array_1509_s104({a_s[1404:0],104'd0},p_prime[104],s_w_104);
AND_array_1509 AND_array_1509_c105({a_c[1403:0],105'd0},p_prime[105],c_w_105);
AND_array_1509 AND_array_1509_s105({a_s[1403:0],105'd0},p_prime[105],s_w_105);
AND_array_1509 AND_array_1509_c106({a_c[1402:0],106'd0},p_prime[106],c_w_106);
AND_array_1509 AND_array_1509_s106({a_s[1402:0],106'd0},p_prime[106],s_w_106);
AND_array_1509 AND_array_1509_c107({a_c[1401:0],107'd0},p_prime[107],c_w_107);
AND_array_1509 AND_array_1509_s107({a_s[1401:0],107'd0},p_prime[107],s_w_107);
AND_array_1509 AND_array_1509_c108({a_c[1400:0],108'd0},p_prime[108],c_w_108);
AND_array_1509 AND_array_1509_s108({a_s[1400:0],108'd0},p_prime[108],s_w_108);
AND_array_1509 AND_array_1509_c109({a_c[1399:0],109'd0},p_prime[109],c_w_109);
AND_array_1509 AND_array_1509_s109({a_s[1399:0],109'd0},p_prime[109],s_w_109);
AND_array_1509 AND_array_1509_c110({a_c[1398:0],110'd0},p_prime[110],c_w_110);
AND_array_1509 AND_array_1509_s110({a_s[1398:0],110'd0},p_prime[110],s_w_110);
AND_array_1509 AND_array_1509_c111({a_c[1397:0],111'd0},p_prime[111],c_w_111);
AND_array_1509 AND_array_1509_s111({a_s[1397:0],111'd0},p_prime[111],s_w_111);
AND_array_1509 AND_array_1509_c112({a_c[1396:0],112'd0},p_prime[112],c_w_112);
AND_array_1509 AND_array_1509_s112({a_s[1396:0],112'd0},p_prime[112],s_w_112);
AND_array_1509 AND_array_1509_c113({a_c[1395:0],113'd0},p_prime[113],c_w_113);
AND_array_1509 AND_array_1509_s113({a_s[1395:0],113'd0},p_prime[113],s_w_113);
AND_array_1509 AND_array_1509_c114({a_c[1394:0],114'd0},p_prime[114],c_w_114);
AND_array_1509 AND_array_1509_s114({a_s[1394:0],114'd0},p_prime[114],s_w_114);
AND_array_1509 AND_array_1509_c115({a_c[1393:0],115'd0},p_prime[115],c_w_115);
AND_array_1509 AND_array_1509_s115({a_s[1393:0],115'd0},p_prime[115],s_w_115);
AND_array_1509 AND_array_1509_c116({a_c[1392:0],116'd0},p_prime[116],c_w_116);
AND_array_1509 AND_array_1509_s116({a_s[1392:0],116'd0},p_prime[116],s_w_116);
AND_array_1509 AND_array_1509_c117({a_c[1391:0],117'd0},p_prime[117],c_w_117);
AND_array_1509 AND_array_1509_s117({a_s[1391:0],117'd0},p_prime[117],s_w_117);
AND_array_1509 AND_array_1509_c118({a_c[1390:0],118'd0},p_prime[118],c_w_118);
AND_array_1509 AND_array_1509_s118({a_s[1390:0],118'd0},p_prime[118],s_w_118);
AND_array_1509 AND_array_1509_c119({a_c[1389:0],119'd0},p_prime[119],c_w_119);
AND_array_1509 AND_array_1509_s119({a_s[1389:0],119'd0},p_prime[119],s_w_119);
AND_array_1509 AND_array_1509_c120({a_c[1388:0],120'd0},p_prime[120],c_w_120);
AND_array_1509 AND_array_1509_s120({a_s[1388:0],120'd0},p_prime[120],s_w_120);
AND_array_1509 AND_array_1509_c121({a_c[1387:0],121'd0},p_prime[121],c_w_121);
AND_array_1509 AND_array_1509_s121({a_s[1387:0],121'd0},p_prime[121],s_w_121);
AND_array_1509 AND_array_1509_c122({a_c[1386:0],122'd0},p_prime[122],c_w_122);
AND_array_1509 AND_array_1509_s122({a_s[1386:0],122'd0},p_prime[122],s_w_122);
AND_array_1509 AND_array_1509_c123({a_c[1385:0],123'd0},p_prime[123],c_w_123);
AND_array_1509 AND_array_1509_s123({a_s[1385:0],123'd0},p_prime[123],s_w_123);
AND_array_1509 AND_array_1509_c124({a_c[1384:0],124'd0},p_prime[124],c_w_124);
AND_array_1509 AND_array_1509_s124({a_s[1384:0],124'd0},p_prime[124],s_w_124);
AND_array_1509 AND_array_1509_c125({a_c[1383:0],125'd0},p_prime[125],c_w_125);
AND_array_1509 AND_array_1509_s125({a_s[1383:0],125'd0},p_prime[125],s_w_125);
AND_array_1509 AND_array_1509_c126({a_c[1382:0],126'd0},p_prime[126],c_w_126);
AND_array_1509 AND_array_1509_s126({a_s[1382:0],126'd0},p_prime[126],s_w_126);
AND_array_1509 AND_array_1509_c127({a_c[1381:0],127'd0},p_prime[127],c_w_127);
AND_array_1509 AND_array_1509_s127({a_s[1381:0],127'd0},p_prime[127],s_w_127);
AND_array_1509 AND_array_1509_c128({a_c[1380:0],128'd0},p_prime[128],c_w_128);
AND_array_1509 AND_array_1509_s128({a_s[1380:0],128'd0},p_prime[128],s_w_128);
AND_array_1509 AND_array_1509_c129({a_c[1379:0],129'd0},p_prime[129],c_w_129);
AND_array_1509 AND_array_1509_s129({a_s[1379:0],129'd0},p_prime[129],s_w_129);
AND_array_1509 AND_array_1509_c130({a_c[1378:0],130'd0},p_prime[130],c_w_130);
AND_array_1509 AND_array_1509_s130({a_s[1378:0],130'd0},p_prime[130],s_w_130);
AND_array_1509 AND_array_1509_c131({a_c[1377:0],131'd0},p_prime[131],c_w_131);
AND_array_1509 AND_array_1509_s131({a_s[1377:0],131'd0},p_prime[131],s_w_131);
AND_array_1509 AND_array_1509_c132({a_c[1376:0],132'd0},p_prime[132],c_w_132);
AND_array_1509 AND_array_1509_s132({a_s[1376:0],132'd0},p_prime[132],s_w_132);
AND_array_1509 AND_array_1509_c133({a_c[1375:0],133'd0},p_prime[133],c_w_133);
AND_array_1509 AND_array_1509_s133({a_s[1375:0],133'd0},p_prime[133],s_w_133);
AND_array_1509 AND_array_1509_c134({a_c[1374:0],134'd0},p_prime[134],c_w_134);
AND_array_1509 AND_array_1509_s134({a_s[1374:0],134'd0},p_prime[134],s_w_134);
AND_array_1509 AND_array_1509_c135({a_c[1373:0],135'd0},p_prime[135],c_w_135);
AND_array_1509 AND_array_1509_s135({a_s[1373:0],135'd0},p_prime[135],s_w_135);
AND_array_1509 AND_array_1509_c136({a_c[1372:0],136'd0},p_prime[136],c_w_136);
AND_array_1509 AND_array_1509_s136({a_s[1372:0],136'd0},p_prime[136],s_w_136);
AND_array_1509 AND_array_1509_c137({a_c[1371:0],137'd0},p_prime[137],c_w_137);
AND_array_1509 AND_array_1509_s137({a_s[1371:0],137'd0},p_prime[137],s_w_137);
AND_array_1509 AND_array_1509_c138({a_c[1370:0],138'd0},p_prime[138],c_w_138);
AND_array_1509 AND_array_1509_s138({a_s[1370:0],138'd0},p_prime[138],s_w_138);
AND_array_1509 AND_array_1509_c139({a_c[1369:0],139'd0},p_prime[139],c_w_139);
AND_array_1509 AND_array_1509_s139({a_s[1369:0],139'd0},p_prime[139],s_w_139);
AND_array_1509 AND_array_1509_c140({a_c[1368:0],140'd0},p_prime[140],c_w_140);
AND_array_1509 AND_array_1509_s140({a_s[1368:0],140'd0},p_prime[140],s_w_140);
AND_array_1509 AND_array_1509_c141({a_c[1367:0],141'd0},p_prime[141],c_w_141);
AND_array_1509 AND_array_1509_s141({a_s[1367:0],141'd0},p_prime[141],s_w_141);
AND_array_1509 AND_array_1509_c142({a_c[1366:0],142'd0},p_prime[142],c_w_142);
AND_array_1509 AND_array_1509_s142({a_s[1366:0],142'd0},p_prime[142],s_w_142);
AND_array_1509 AND_array_1509_c143({a_c[1365:0],143'd0},p_prime[143],c_w_143);
AND_array_1509 AND_array_1509_s143({a_s[1365:0],143'd0},p_prime[143],s_w_143);
AND_array_1509 AND_array_1509_c144({a_c[1364:0],144'd0},p_prime[144],c_w_144);
AND_array_1509 AND_array_1509_s144({a_s[1364:0],144'd0},p_prime[144],s_w_144);
AND_array_1509 AND_array_1509_c145({a_c[1363:0],145'd0},p_prime[145],c_w_145);
AND_array_1509 AND_array_1509_s145({a_s[1363:0],145'd0},p_prime[145],s_w_145);
AND_array_1509 AND_array_1509_c146({a_c[1362:0],146'd0},p_prime[146],c_w_146);
AND_array_1509 AND_array_1509_s146({a_s[1362:0],146'd0},p_prime[146],s_w_146);
AND_array_1509 AND_array_1509_c147({a_c[1361:0],147'd0},p_prime[147],c_w_147);
AND_array_1509 AND_array_1509_s147({a_s[1361:0],147'd0},p_prime[147],s_w_147);
AND_array_1509 AND_array_1509_c148({a_c[1360:0],148'd0},p_prime[148],c_w_148);
AND_array_1509 AND_array_1509_s148({a_s[1360:0],148'd0},p_prime[148],s_w_148);
AND_array_1509 AND_array_1509_c149({a_c[1359:0],149'd0},p_prime[149],c_w_149);
AND_array_1509 AND_array_1509_s149({a_s[1359:0],149'd0},p_prime[149],s_w_149);
AND_array_1509 AND_array_1509_c150({a_c[1358:0],150'd0},p_prime[150],c_w_150);
AND_array_1509 AND_array_1509_s150({a_s[1358:0],150'd0},p_prime[150],s_w_150);
AND_array_1509 AND_array_1509_c151({a_c[1357:0],151'd0},p_prime[151],c_w_151);
AND_array_1509 AND_array_1509_s151({a_s[1357:0],151'd0},p_prime[151],s_w_151);
AND_array_1509 AND_array_1509_c152({a_c[1356:0],152'd0},p_prime[152],c_w_152);
AND_array_1509 AND_array_1509_s152({a_s[1356:0],152'd0},p_prime[152],s_w_152);
AND_array_1509 AND_array_1509_c153({a_c[1355:0],153'd0},p_prime[153],c_w_153);
AND_array_1509 AND_array_1509_s153({a_s[1355:0],153'd0},p_prime[153],s_w_153);
AND_array_1509 AND_array_1509_c154({a_c[1354:0],154'd0},p_prime[154],c_w_154);
AND_array_1509 AND_array_1509_s154({a_s[1354:0],154'd0},p_prime[154],s_w_154);
AND_array_1509 AND_array_1509_c155({a_c[1353:0],155'd0},p_prime[155],c_w_155);
AND_array_1509 AND_array_1509_s155({a_s[1353:0],155'd0},p_prime[155],s_w_155);
AND_array_1509 AND_array_1509_c156({a_c[1352:0],156'd0},p_prime[156],c_w_156);
AND_array_1509 AND_array_1509_s156({a_s[1352:0],156'd0},p_prime[156],s_w_156);
AND_array_1509 AND_array_1509_c157({a_c[1351:0],157'd0},p_prime[157],c_w_157);
AND_array_1509 AND_array_1509_s157({a_s[1351:0],157'd0},p_prime[157],s_w_157);
AND_array_1509 AND_array_1509_c158({a_c[1350:0],158'd0},p_prime[158],c_w_158);
AND_array_1509 AND_array_1509_s158({a_s[1350:0],158'd0},p_prime[158],s_w_158);
AND_array_1509 AND_array_1509_c159({a_c[1349:0],159'd0},p_prime[159],c_w_159);
AND_array_1509 AND_array_1509_s159({a_s[1349:0],159'd0},p_prime[159],s_w_159);
AND_array_1509 AND_array_1509_c160({a_c[1348:0],160'd0},p_prime[160],c_w_160);
AND_array_1509 AND_array_1509_s160({a_s[1348:0],160'd0},p_prime[160],s_w_160);
AND_array_1509 AND_array_1509_c161({a_c[1347:0],161'd0},p_prime[161],c_w_161);
AND_array_1509 AND_array_1509_s161({a_s[1347:0],161'd0},p_prime[161],s_w_161);
AND_array_1509 AND_array_1509_c162({a_c[1346:0],162'd0},p_prime[162],c_w_162);
AND_array_1509 AND_array_1509_s162({a_s[1346:0],162'd0},p_prime[162],s_w_162);
AND_array_1509 AND_array_1509_c163({a_c[1345:0],163'd0},p_prime[163],c_w_163);
AND_array_1509 AND_array_1509_s163({a_s[1345:0],163'd0},p_prime[163],s_w_163);
AND_array_1509 AND_array_1509_c164({a_c[1344:0],164'd0},p_prime[164],c_w_164);
AND_array_1509 AND_array_1509_s164({a_s[1344:0],164'd0},p_prime[164],s_w_164);
AND_array_1509 AND_array_1509_c165({a_c[1343:0],165'd0},p_prime[165],c_w_165);
AND_array_1509 AND_array_1509_s165({a_s[1343:0],165'd0},p_prime[165],s_w_165);
AND_array_1509 AND_array_1509_c166({a_c[1342:0],166'd0},p_prime[166],c_w_166);
AND_array_1509 AND_array_1509_s166({a_s[1342:0],166'd0},p_prime[166],s_w_166);
AND_array_1509 AND_array_1509_c167({a_c[1341:0],167'd0},p_prime[167],c_w_167);
AND_array_1509 AND_array_1509_s167({a_s[1341:0],167'd0},p_prime[167],s_w_167);
AND_array_1509 AND_array_1509_c168({a_c[1340:0],168'd0},p_prime[168],c_w_168);
AND_array_1509 AND_array_1509_s168({a_s[1340:0],168'd0},p_prime[168],s_w_168);
AND_array_1509 AND_array_1509_c169({a_c[1339:0],169'd0},p_prime[169],c_w_169);
AND_array_1509 AND_array_1509_s169({a_s[1339:0],169'd0},p_prime[169],s_w_169);
AND_array_1509 AND_array_1509_c170({a_c[1338:0],170'd0},p_prime[170],c_w_170);
AND_array_1509 AND_array_1509_s170({a_s[1338:0],170'd0},p_prime[170],s_w_170);
AND_array_1509 AND_array_1509_c171({a_c[1337:0],171'd0},p_prime[171],c_w_171);
AND_array_1509 AND_array_1509_s171({a_s[1337:0],171'd0},p_prime[171],s_w_171);
AND_array_1509 AND_array_1509_c172({a_c[1336:0],172'd0},p_prime[172],c_w_172);
AND_array_1509 AND_array_1509_s172({a_s[1336:0],172'd0},p_prime[172],s_w_172);
AND_array_1509 AND_array_1509_c173({a_c[1335:0],173'd0},p_prime[173],c_w_173);
AND_array_1509 AND_array_1509_s173({a_s[1335:0],173'd0},p_prime[173],s_w_173);
AND_array_1509 AND_array_1509_c174({a_c[1334:0],174'd0},p_prime[174],c_w_174);
AND_array_1509 AND_array_1509_s174({a_s[1334:0],174'd0},p_prime[174],s_w_174);
AND_array_1509 AND_array_1509_c175({a_c[1333:0],175'd0},p_prime[175],c_w_175);
AND_array_1509 AND_array_1509_s175({a_s[1333:0],175'd0},p_prime[175],s_w_175);
AND_array_1509 AND_array_1509_c176({a_c[1332:0],176'd0},p_prime[176],c_w_176);
AND_array_1509 AND_array_1509_s176({a_s[1332:0],176'd0},p_prime[176],s_w_176);
AND_array_1509 AND_array_1509_c177({a_c[1331:0],177'd0},p_prime[177],c_w_177);
AND_array_1509 AND_array_1509_s177({a_s[1331:0],177'd0},p_prime[177],s_w_177);
AND_array_1509 AND_array_1509_c178({a_c[1330:0],178'd0},p_prime[178],c_w_178);
AND_array_1509 AND_array_1509_s178({a_s[1330:0],178'd0},p_prime[178],s_w_178);
AND_array_1509 AND_array_1509_c179({a_c[1329:0],179'd0},p_prime[179],c_w_179);
AND_array_1509 AND_array_1509_s179({a_s[1329:0],179'd0},p_prime[179],s_w_179);
AND_array_1509 AND_array_1509_c180({a_c[1328:0],180'd0},p_prime[180],c_w_180);
AND_array_1509 AND_array_1509_s180({a_s[1328:0],180'd0},p_prime[180],s_w_180);
AND_array_1509 AND_array_1509_c181({a_c[1327:0],181'd0},p_prime[181],c_w_181);
AND_array_1509 AND_array_1509_s181({a_s[1327:0],181'd0},p_prime[181],s_w_181);
AND_array_1509 AND_array_1509_c182({a_c[1326:0],182'd0},p_prime[182],c_w_182);
AND_array_1509 AND_array_1509_s182({a_s[1326:0],182'd0},p_prime[182],s_w_182);
AND_array_1509 AND_array_1509_c183({a_c[1325:0],183'd0},p_prime[183],c_w_183);
AND_array_1509 AND_array_1509_s183({a_s[1325:0],183'd0},p_prime[183],s_w_183);
AND_array_1509 AND_array_1509_c184({a_c[1324:0],184'd0},p_prime[184],c_w_184);
AND_array_1509 AND_array_1509_s184({a_s[1324:0],184'd0},p_prime[184],s_w_184);
AND_array_1509 AND_array_1509_c185({a_c[1323:0],185'd0},p_prime[185],c_w_185);
AND_array_1509 AND_array_1509_s185({a_s[1323:0],185'd0},p_prime[185],s_w_185);
AND_array_1509 AND_array_1509_c186({a_c[1322:0],186'd0},p_prime[186],c_w_186);
AND_array_1509 AND_array_1509_s186({a_s[1322:0],186'd0},p_prime[186],s_w_186);
AND_array_1509 AND_array_1509_c187({a_c[1321:0],187'd0},p_prime[187],c_w_187);
AND_array_1509 AND_array_1509_s187({a_s[1321:0],187'd0},p_prime[187],s_w_187);
AND_array_1509 AND_array_1509_c188({a_c[1320:0],188'd0},p_prime[188],c_w_188);
AND_array_1509 AND_array_1509_s188({a_s[1320:0],188'd0},p_prime[188],s_w_188);
AND_array_1509 AND_array_1509_c189({a_c[1319:0],189'd0},p_prime[189],c_w_189);
AND_array_1509 AND_array_1509_s189({a_s[1319:0],189'd0},p_prime[189],s_w_189);
AND_array_1509 AND_array_1509_c190({a_c[1318:0],190'd0},p_prime[190],c_w_190);
AND_array_1509 AND_array_1509_s190({a_s[1318:0],190'd0},p_prime[190],s_w_190);
AND_array_1509 AND_array_1509_c191({a_c[1317:0],191'd0},p_prime[191],c_w_191);
AND_array_1509 AND_array_1509_s191({a_s[1317:0],191'd0},p_prime[191],s_w_191);
AND_array_1509 AND_array_1509_c192({a_c[1316:0],192'd0},p_prime[192],c_w_192);
AND_array_1509 AND_array_1509_s192({a_s[1316:0],192'd0},p_prime[192],s_w_192);
AND_array_1509 AND_array_1509_c193({a_c[1315:0],193'd0},p_prime[193],c_w_193);
AND_array_1509 AND_array_1509_s193({a_s[1315:0],193'd0},p_prime[193],s_w_193);
AND_array_1509 AND_array_1509_c194({a_c[1314:0],194'd0},p_prime[194],c_w_194);
AND_array_1509 AND_array_1509_s194({a_s[1314:0],194'd0},p_prime[194],s_w_194);
AND_array_1509 AND_array_1509_c195({a_c[1313:0],195'd0},p_prime[195],c_w_195);
AND_array_1509 AND_array_1509_s195({a_s[1313:0],195'd0},p_prime[195],s_w_195);
AND_array_1509 AND_array_1509_c196({a_c[1312:0],196'd0},p_prime[196],c_w_196);
AND_array_1509 AND_array_1509_s196({a_s[1312:0],196'd0},p_prime[196],s_w_196);
AND_array_1509 AND_array_1509_c197({a_c[1311:0],197'd0},p_prime[197],c_w_197);
AND_array_1509 AND_array_1509_s197({a_s[1311:0],197'd0},p_prime[197],s_w_197);
AND_array_1509 AND_array_1509_c198({a_c[1310:0],198'd0},p_prime[198],c_w_198);
AND_array_1509 AND_array_1509_s198({a_s[1310:0],198'd0},p_prime[198],s_w_198);
AND_array_1509 AND_array_1509_c199({a_c[1309:0],199'd0},p_prime[199],c_w_199);
AND_array_1509 AND_array_1509_s199({a_s[1309:0],199'd0},p_prime[199],s_w_199);
AND_array_1509 AND_array_1509_c200({a_c[1308:0],200'd0},p_prime[200],c_w_200);
AND_array_1509 AND_array_1509_s200({a_s[1308:0],200'd0},p_prime[200],s_w_200);
AND_array_1509 AND_array_1509_c201({a_c[1307:0],201'd0},p_prime[201],c_w_201);
AND_array_1509 AND_array_1509_s201({a_s[1307:0],201'd0},p_prime[201],s_w_201);
AND_array_1509 AND_array_1509_c202({a_c[1306:0],202'd0},p_prime[202],c_w_202);
AND_array_1509 AND_array_1509_s202({a_s[1306:0],202'd0},p_prime[202],s_w_202);
AND_array_1509 AND_array_1509_c203({a_c[1305:0],203'd0},p_prime[203],c_w_203);
AND_array_1509 AND_array_1509_s203({a_s[1305:0],203'd0},p_prime[203],s_w_203);
AND_array_1509 AND_array_1509_c204({a_c[1304:0],204'd0},p_prime[204],c_w_204);
AND_array_1509 AND_array_1509_s204({a_s[1304:0],204'd0},p_prime[204],s_w_204);
AND_array_1509 AND_array_1509_c205({a_c[1303:0],205'd0},p_prime[205],c_w_205);
AND_array_1509 AND_array_1509_s205({a_s[1303:0],205'd0},p_prime[205],s_w_205);
AND_array_1509 AND_array_1509_c206({a_c[1302:0],206'd0},p_prime[206],c_w_206);
AND_array_1509 AND_array_1509_s206({a_s[1302:0],206'd0},p_prime[206],s_w_206);
AND_array_1509 AND_array_1509_c207({a_c[1301:0],207'd0},p_prime[207],c_w_207);
AND_array_1509 AND_array_1509_s207({a_s[1301:0],207'd0},p_prime[207],s_w_207);
AND_array_1509 AND_array_1509_c208({a_c[1300:0],208'd0},p_prime[208],c_w_208);
AND_array_1509 AND_array_1509_s208({a_s[1300:0],208'd0},p_prime[208],s_w_208);
AND_array_1509 AND_array_1509_c209({a_c[1299:0],209'd0},p_prime[209],c_w_209);
AND_array_1509 AND_array_1509_s209({a_s[1299:0],209'd0},p_prime[209],s_w_209);
AND_array_1509 AND_array_1509_c210({a_c[1298:0],210'd0},p_prime[210],c_w_210);
AND_array_1509 AND_array_1509_s210({a_s[1298:0],210'd0},p_prime[210],s_w_210);
AND_array_1509 AND_array_1509_c211({a_c[1297:0],211'd0},p_prime[211],c_w_211);
AND_array_1509 AND_array_1509_s211({a_s[1297:0],211'd0},p_prime[211],s_w_211);
AND_array_1509 AND_array_1509_c212({a_c[1296:0],212'd0},p_prime[212],c_w_212);
AND_array_1509 AND_array_1509_s212({a_s[1296:0],212'd0},p_prime[212],s_w_212);
AND_array_1509 AND_array_1509_c213({a_c[1295:0],213'd0},p_prime[213],c_w_213);
AND_array_1509 AND_array_1509_s213({a_s[1295:0],213'd0},p_prime[213],s_w_213);
AND_array_1509 AND_array_1509_c214({a_c[1294:0],214'd0},p_prime[214],c_w_214);
AND_array_1509 AND_array_1509_s214({a_s[1294:0],214'd0},p_prime[214],s_w_214);
AND_array_1509 AND_array_1509_c215({a_c[1293:0],215'd0},p_prime[215],c_w_215);
AND_array_1509 AND_array_1509_s215({a_s[1293:0],215'd0},p_prime[215],s_w_215);
AND_array_1509 AND_array_1509_c216({a_c[1292:0],216'd0},p_prime[216],c_w_216);
AND_array_1509 AND_array_1509_s216({a_s[1292:0],216'd0},p_prime[216],s_w_216);
AND_array_1509 AND_array_1509_c217({a_c[1291:0],217'd0},p_prime[217],c_w_217);
AND_array_1509 AND_array_1509_s217({a_s[1291:0],217'd0},p_prime[217],s_w_217);
AND_array_1509 AND_array_1509_c218({a_c[1290:0],218'd0},p_prime[218],c_w_218);
AND_array_1509 AND_array_1509_s218({a_s[1290:0],218'd0},p_prime[218],s_w_218);
AND_array_1509 AND_array_1509_c219({a_c[1289:0],219'd0},p_prime[219],c_w_219);
AND_array_1509 AND_array_1509_s219({a_s[1289:0],219'd0},p_prime[219],s_w_219);
AND_array_1509 AND_array_1509_c220({a_c[1288:0],220'd0},p_prime[220],c_w_220);
AND_array_1509 AND_array_1509_s220({a_s[1288:0],220'd0},p_prime[220],s_w_220);
AND_array_1509 AND_array_1509_c221({a_c[1287:0],221'd0},p_prime[221],c_w_221);
AND_array_1509 AND_array_1509_s221({a_s[1287:0],221'd0},p_prime[221],s_w_221);
AND_array_1509 AND_array_1509_c222({a_c[1286:0],222'd0},p_prime[222],c_w_222);
AND_array_1509 AND_array_1509_s222({a_s[1286:0],222'd0},p_prime[222],s_w_222);
AND_array_1509 AND_array_1509_c223({a_c[1285:0],223'd0},p_prime[223],c_w_223);
AND_array_1509 AND_array_1509_s223({a_s[1285:0],223'd0},p_prime[223],s_w_223);
AND_array_1509 AND_array_1509_c224({a_c[1284:0],224'd0},p_prime[224],c_w_224);
AND_array_1509 AND_array_1509_s224({a_s[1284:0],224'd0},p_prime[224],s_w_224);
AND_array_1509 AND_array_1509_c225({a_c[1283:0],225'd0},p_prime[225],c_w_225);
AND_array_1509 AND_array_1509_s225({a_s[1283:0],225'd0},p_prime[225],s_w_225);
AND_array_1509 AND_array_1509_c226({a_c[1282:0],226'd0},p_prime[226],c_w_226);
AND_array_1509 AND_array_1509_s226({a_s[1282:0],226'd0},p_prime[226],s_w_226);
AND_array_1509 AND_array_1509_c227({a_c[1281:0],227'd0},p_prime[227],c_w_227);
AND_array_1509 AND_array_1509_s227({a_s[1281:0],227'd0},p_prime[227],s_w_227);
AND_array_1509 AND_array_1509_c228({a_c[1280:0],228'd0},p_prime[228],c_w_228);
AND_array_1509 AND_array_1509_s228({a_s[1280:0],228'd0},p_prime[228],s_w_228);
AND_array_1509 AND_array_1509_c229({a_c[1279:0],229'd0},p_prime[229],c_w_229);
AND_array_1509 AND_array_1509_s229({a_s[1279:0],229'd0},p_prime[229],s_w_229);
AND_array_1509 AND_array_1509_c230({a_c[1278:0],230'd0},p_prime[230],c_w_230);
AND_array_1509 AND_array_1509_s230({a_s[1278:0],230'd0},p_prime[230],s_w_230);
AND_array_1509 AND_array_1509_c231({a_c[1277:0],231'd0},p_prime[231],c_w_231);
AND_array_1509 AND_array_1509_s231({a_s[1277:0],231'd0},p_prime[231],s_w_231);
AND_array_1509 AND_array_1509_c232({a_c[1276:0],232'd0},p_prime[232],c_w_232);
AND_array_1509 AND_array_1509_s232({a_s[1276:0],232'd0},p_prime[232],s_w_232);
AND_array_1509 AND_array_1509_c233({a_c[1275:0],233'd0},p_prime[233],c_w_233);
AND_array_1509 AND_array_1509_s233({a_s[1275:0],233'd0},p_prime[233],s_w_233);
AND_array_1509 AND_array_1509_c234({a_c[1274:0],234'd0},p_prime[234],c_w_234);
AND_array_1509 AND_array_1509_s234({a_s[1274:0],234'd0},p_prime[234],s_w_234);
AND_array_1509 AND_array_1509_c235({a_c[1273:0],235'd0},p_prime[235],c_w_235);
AND_array_1509 AND_array_1509_s235({a_s[1273:0],235'd0},p_prime[235],s_w_235);
AND_array_1509 AND_array_1509_c236({a_c[1272:0],236'd0},p_prime[236],c_w_236);
AND_array_1509 AND_array_1509_s236({a_s[1272:0],236'd0},p_prime[236],s_w_236);
AND_array_1509 AND_array_1509_c237({a_c[1271:0],237'd0},p_prime[237],c_w_237);
AND_array_1509 AND_array_1509_s237({a_s[1271:0],237'd0},p_prime[237],s_w_237);
AND_array_1509 AND_array_1509_c238({a_c[1270:0],238'd0},p_prime[238],c_w_238);
AND_array_1509 AND_array_1509_s238({a_s[1270:0],238'd0},p_prime[238],s_w_238);
AND_array_1509 AND_array_1509_c239({a_c[1269:0],239'd0},p_prime[239],c_w_239);
AND_array_1509 AND_array_1509_s239({a_s[1269:0],239'd0},p_prime[239],s_w_239);
AND_array_1509 AND_array_1509_c240({a_c[1268:0],240'd0},p_prime[240],c_w_240);
AND_array_1509 AND_array_1509_s240({a_s[1268:0],240'd0},p_prime[240],s_w_240);
AND_array_1509 AND_array_1509_c241({a_c[1267:0],241'd0},p_prime[241],c_w_241);
AND_array_1509 AND_array_1509_s241({a_s[1267:0],241'd0},p_prime[241],s_w_241);
AND_array_1509 AND_array_1509_c242({a_c[1266:0],242'd0},p_prime[242],c_w_242);
AND_array_1509 AND_array_1509_s242({a_s[1266:0],242'd0},p_prime[242],s_w_242);
AND_array_1509 AND_array_1509_c243({a_c[1265:0],243'd0},p_prime[243],c_w_243);
AND_array_1509 AND_array_1509_s243({a_s[1265:0],243'd0},p_prime[243],s_w_243);
AND_array_1509 AND_array_1509_c244({a_c[1264:0],244'd0},p_prime[244],c_w_244);
AND_array_1509 AND_array_1509_s244({a_s[1264:0],244'd0},p_prime[244],s_w_244);
AND_array_1509 AND_array_1509_c245({a_c[1263:0],245'd0},p_prime[245],c_w_245);
AND_array_1509 AND_array_1509_s245({a_s[1263:0],245'd0},p_prime[245],s_w_245);
AND_array_1509 AND_array_1509_c246({a_c[1262:0],246'd0},p_prime[246],c_w_246);
AND_array_1509 AND_array_1509_s246({a_s[1262:0],246'd0},p_prime[246],s_w_246);
AND_array_1509 AND_array_1509_c247({a_c[1261:0],247'd0},p_prime[247],c_w_247);
AND_array_1509 AND_array_1509_s247({a_s[1261:0],247'd0},p_prime[247],s_w_247);
AND_array_1509 AND_array_1509_c248({a_c[1260:0],248'd0},p_prime[248],c_w_248);
AND_array_1509 AND_array_1509_s248({a_s[1260:0],248'd0},p_prime[248],s_w_248);
AND_array_1509 AND_array_1509_c249({a_c[1259:0],249'd0},p_prime[249],c_w_249);
AND_array_1509 AND_array_1509_s249({a_s[1259:0],249'd0},p_prime[249],s_w_249);
AND_array_1509 AND_array_1509_c250({a_c[1258:0],250'd0},p_prime[250],c_w_250);
AND_array_1509 AND_array_1509_s250({a_s[1258:0],250'd0},p_prime[250],s_w_250);
AND_array_1509 AND_array_1509_c251({a_c[1257:0],251'd0},p_prime[251],c_w_251);
AND_array_1509 AND_array_1509_s251({a_s[1257:0],251'd0},p_prime[251],s_w_251);
AND_array_1509 AND_array_1509_c252({a_c[1256:0],252'd0},p_prime[252],c_w_252);
AND_array_1509 AND_array_1509_s252({a_s[1256:0],252'd0},p_prime[252],s_w_252);
AND_array_1509 AND_array_1509_c253({a_c[1255:0],253'd0},p_prime[253],c_w_253);
AND_array_1509 AND_array_1509_s253({a_s[1255:0],253'd0},p_prime[253],s_w_253);
AND_array_1509 AND_array_1509_c254({a_c[1254:0],254'd0},p_prime[254],c_w_254);
AND_array_1509 AND_array_1509_s254({a_s[1254:0],254'd0},p_prime[254],s_w_254);
AND_array_1509 AND_array_1509_c255({a_c[1253:0],255'd0},p_prime[255],c_w_255);
AND_array_1509 AND_array_1509_s255({a_s[1253:0],255'd0},p_prime[255],s_w_255);
AND_array_1509 AND_array_1509_c256({a_c[1252:0],256'd0},p_prime[256],c_w_256);
AND_array_1509 AND_array_1509_s256({a_s[1252:0],256'd0},p_prime[256],s_w_256);
AND_array_1509 AND_array_1509_c257({a_c[1251:0],257'd0},p_prime[257],c_w_257);
AND_array_1509 AND_array_1509_s257({a_s[1251:0],257'd0},p_prime[257],s_w_257);
AND_array_1509 AND_array_1509_c258({a_c[1250:0],258'd0},p_prime[258],c_w_258);
AND_array_1509 AND_array_1509_s258({a_s[1250:0],258'd0},p_prime[258],s_w_258);
AND_array_1509 AND_array_1509_c259({a_c[1249:0],259'd0},p_prime[259],c_w_259);
AND_array_1509 AND_array_1509_s259({a_s[1249:0],259'd0},p_prime[259],s_w_259);
AND_array_1509 AND_array_1509_c260({a_c[1248:0],260'd0},p_prime[260],c_w_260);
AND_array_1509 AND_array_1509_s260({a_s[1248:0],260'd0},p_prime[260],s_w_260);
AND_array_1509 AND_array_1509_c261({a_c[1247:0],261'd0},p_prime[261],c_w_261);
AND_array_1509 AND_array_1509_s261({a_s[1247:0],261'd0},p_prime[261],s_w_261);
AND_array_1509 AND_array_1509_c262({a_c[1246:0],262'd0},p_prime[262],c_w_262);
AND_array_1509 AND_array_1509_s262({a_s[1246:0],262'd0},p_prime[262],s_w_262);
AND_array_1509 AND_array_1509_c263({a_c[1245:0],263'd0},p_prime[263],c_w_263);
AND_array_1509 AND_array_1509_s263({a_s[1245:0],263'd0},p_prime[263],s_w_263);
AND_array_1509 AND_array_1509_c264({a_c[1244:0],264'd0},p_prime[264],c_w_264);
AND_array_1509 AND_array_1509_s264({a_s[1244:0],264'd0},p_prime[264],s_w_264);
AND_array_1509 AND_array_1509_c265({a_c[1243:0],265'd0},p_prime[265],c_w_265);
AND_array_1509 AND_array_1509_s265({a_s[1243:0],265'd0},p_prime[265],s_w_265);
AND_array_1509 AND_array_1509_c266({a_c[1242:0],266'd0},p_prime[266],c_w_266);
AND_array_1509 AND_array_1509_s266({a_s[1242:0],266'd0},p_prime[266],s_w_266);
AND_array_1509 AND_array_1509_c267({a_c[1241:0],267'd0},p_prime[267],c_w_267);
AND_array_1509 AND_array_1509_s267({a_s[1241:0],267'd0},p_prime[267],s_w_267);
AND_array_1509 AND_array_1509_c268({a_c[1240:0],268'd0},p_prime[268],c_w_268);
AND_array_1509 AND_array_1509_s268({a_s[1240:0],268'd0},p_prime[268],s_w_268);
AND_array_1509 AND_array_1509_c269({a_c[1239:0],269'd0},p_prime[269],c_w_269);
AND_array_1509 AND_array_1509_s269({a_s[1239:0],269'd0},p_prime[269],s_w_269);
AND_array_1509 AND_array_1509_c270({a_c[1238:0],270'd0},p_prime[270],c_w_270);
AND_array_1509 AND_array_1509_s270({a_s[1238:0],270'd0},p_prime[270],s_w_270);
AND_array_1509 AND_array_1509_c271({a_c[1237:0],271'd0},p_prime[271],c_w_271);
AND_array_1509 AND_array_1509_s271({a_s[1237:0],271'd0},p_prime[271],s_w_271);
AND_array_1509 AND_array_1509_c272({a_c[1236:0],272'd0},p_prime[272],c_w_272);
AND_array_1509 AND_array_1509_s272({a_s[1236:0],272'd0},p_prime[272],s_w_272);
AND_array_1509 AND_array_1509_c273({a_c[1235:0],273'd0},p_prime[273],c_w_273);
AND_array_1509 AND_array_1509_s273({a_s[1235:0],273'd0},p_prime[273],s_w_273);
AND_array_1509 AND_array_1509_c274({a_c[1234:0],274'd0},p_prime[274],c_w_274);
AND_array_1509 AND_array_1509_s274({a_s[1234:0],274'd0},p_prime[274],s_w_274);
AND_array_1509 AND_array_1509_c275({a_c[1233:0],275'd0},p_prime[275],c_w_275);
AND_array_1509 AND_array_1509_s275({a_s[1233:0],275'd0},p_prime[275],s_w_275);
AND_array_1509 AND_array_1509_c276({a_c[1232:0],276'd0},p_prime[276],c_w_276);
AND_array_1509 AND_array_1509_s276({a_s[1232:0],276'd0},p_prime[276],s_w_276);
AND_array_1509 AND_array_1509_c277({a_c[1231:0],277'd0},p_prime[277],c_w_277);
AND_array_1509 AND_array_1509_s277({a_s[1231:0],277'd0},p_prime[277],s_w_277);
AND_array_1509 AND_array_1509_c278({a_c[1230:0],278'd0},p_prime[278],c_w_278);
AND_array_1509 AND_array_1509_s278({a_s[1230:0],278'd0},p_prime[278],s_w_278);
AND_array_1509 AND_array_1509_c279({a_c[1229:0],279'd0},p_prime[279],c_w_279);
AND_array_1509 AND_array_1509_s279({a_s[1229:0],279'd0},p_prime[279],s_w_279);
AND_array_1509 AND_array_1509_c280({a_c[1228:0],280'd0},p_prime[280],c_w_280);
AND_array_1509 AND_array_1509_s280({a_s[1228:0],280'd0},p_prime[280],s_w_280);
AND_array_1509 AND_array_1509_c281({a_c[1227:0],281'd0},p_prime[281],c_w_281);
AND_array_1509 AND_array_1509_s281({a_s[1227:0],281'd0},p_prime[281],s_w_281);
AND_array_1509 AND_array_1509_c282({a_c[1226:0],282'd0},p_prime[282],c_w_282);
AND_array_1509 AND_array_1509_s282({a_s[1226:0],282'd0},p_prime[282],s_w_282);
AND_array_1509 AND_array_1509_c283({a_c[1225:0],283'd0},p_prime[283],c_w_283);
AND_array_1509 AND_array_1509_s283({a_s[1225:0],283'd0},p_prime[283],s_w_283);
AND_array_1509 AND_array_1509_c284({a_c[1224:0],284'd0},p_prime[284],c_w_284);
AND_array_1509 AND_array_1509_s284({a_s[1224:0],284'd0},p_prime[284],s_w_284);
AND_array_1509 AND_array_1509_c285({a_c[1223:0],285'd0},p_prime[285],c_w_285);
AND_array_1509 AND_array_1509_s285({a_s[1223:0],285'd0},p_prime[285],s_w_285);
AND_array_1509 AND_array_1509_c286({a_c[1222:0],286'd0},p_prime[286],c_w_286);
AND_array_1509 AND_array_1509_s286({a_s[1222:0],286'd0},p_prime[286],s_w_286);
AND_array_1509 AND_array_1509_c287({a_c[1221:0],287'd0},p_prime[287],c_w_287);
AND_array_1509 AND_array_1509_s287({a_s[1221:0],287'd0},p_prime[287],s_w_287);
AND_array_1509 AND_array_1509_c288({a_c[1220:0],288'd0},p_prime[288],c_w_288);
AND_array_1509 AND_array_1509_s288({a_s[1220:0],288'd0},p_prime[288],s_w_288);
AND_array_1509 AND_array_1509_c289({a_c[1219:0],289'd0},p_prime[289],c_w_289);
AND_array_1509 AND_array_1509_s289({a_s[1219:0],289'd0},p_prime[289],s_w_289);
AND_array_1509 AND_array_1509_c290({a_c[1218:0],290'd0},p_prime[290],c_w_290);
AND_array_1509 AND_array_1509_s290({a_s[1218:0],290'd0},p_prime[290],s_w_290);
AND_array_1509 AND_array_1509_c291({a_c[1217:0],291'd0},p_prime[291],c_w_291);
AND_array_1509 AND_array_1509_s291({a_s[1217:0],291'd0},p_prime[291],s_w_291);
AND_array_1509 AND_array_1509_c292({a_c[1216:0],292'd0},p_prime[292],c_w_292);
AND_array_1509 AND_array_1509_s292({a_s[1216:0],292'd0},p_prime[292],s_w_292);
AND_array_1509 AND_array_1509_c293({a_c[1215:0],293'd0},p_prime[293],c_w_293);
AND_array_1509 AND_array_1509_s293({a_s[1215:0],293'd0},p_prime[293],s_w_293);
AND_array_1509 AND_array_1509_c294({a_c[1214:0],294'd0},p_prime[294],c_w_294);
AND_array_1509 AND_array_1509_s294({a_s[1214:0],294'd0},p_prime[294],s_w_294);
AND_array_1509 AND_array_1509_c295({a_c[1213:0],295'd0},p_prime[295],c_w_295);
AND_array_1509 AND_array_1509_s295({a_s[1213:0],295'd0},p_prime[295],s_w_295);
AND_array_1509 AND_array_1509_c296({a_c[1212:0],296'd0},p_prime[296],c_w_296);
AND_array_1509 AND_array_1509_s296({a_s[1212:0],296'd0},p_prime[296],s_w_296);
AND_array_1509 AND_array_1509_c297({a_c[1211:0],297'd0},p_prime[297],c_w_297);
AND_array_1509 AND_array_1509_s297({a_s[1211:0],297'd0},p_prime[297],s_w_297);
AND_array_1509 AND_array_1509_c298({a_c[1210:0],298'd0},p_prime[298],c_w_298);
AND_array_1509 AND_array_1509_s298({a_s[1210:0],298'd0},p_prime[298],s_w_298);
AND_array_1509 AND_array_1509_c299({a_c[1209:0],299'd0},p_prime[299],c_w_299);
AND_array_1509 AND_array_1509_s299({a_s[1209:0],299'd0},p_prime[299],s_w_299);
AND_array_1509 AND_array_1509_c300({a_c[1208:0],300'd0},p_prime[300],c_w_300);
AND_array_1509 AND_array_1509_s300({a_s[1208:0],300'd0},p_prime[300],s_w_300);
AND_array_1509 AND_array_1509_c301({a_c[1207:0],301'd0},p_prime[301],c_w_301);
AND_array_1509 AND_array_1509_s301({a_s[1207:0],301'd0},p_prime[301],s_w_301);
AND_array_1509 AND_array_1509_c302({a_c[1206:0],302'd0},p_prime[302],c_w_302);
AND_array_1509 AND_array_1509_s302({a_s[1206:0],302'd0},p_prime[302],s_w_302);
AND_array_1509 AND_array_1509_c303({a_c[1205:0],303'd0},p_prime[303],c_w_303);
AND_array_1509 AND_array_1509_s303({a_s[1205:0],303'd0},p_prime[303],s_w_303);
AND_array_1509 AND_array_1509_c304({a_c[1204:0],304'd0},p_prime[304],c_w_304);
AND_array_1509 AND_array_1509_s304({a_s[1204:0],304'd0},p_prime[304],s_w_304);
AND_array_1509 AND_array_1509_c305({a_c[1203:0],305'd0},p_prime[305],c_w_305);
AND_array_1509 AND_array_1509_s305({a_s[1203:0],305'd0},p_prime[305],s_w_305);
AND_array_1509 AND_array_1509_c306({a_c[1202:0],306'd0},p_prime[306],c_w_306);
AND_array_1509 AND_array_1509_s306({a_s[1202:0],306'd0},p_prime[306],s_w_306);
AND_array_1509 AND_array_1509_c307({a_c[1201:0],307'd0},p_prime[307],c_w_307);
AND_array_1509 AND_array_1509_s307({a_s[1201:0],307'd0},p_prime[307],s_w_307);
AND_array_1509 AND_array_1509_c308({a_c[1200:0],308'd0},p_prime[308],c_w_308);
AND_array_1509 AND_array_1509_s308({a_s[1200:0],308'd0},p_prime[308],s_w_308);
AND_array_1509 AND_array_1509_c309({a_c[1199:0],309'd0},p_prime[309],c_w_309);
AND_array_1509 AND_array_1509_s309({a_s[1199:0],309'd0},p_prime[309],s_w_309);
AND_array_1509 AND_array_1509_c310({a_c[1198:0],310'd0},p_prime[310],c_w_310);
AND_array_1509 AND_array_1509_s310({a_s[1198:0],310'd0},p_prime[310],s_w_310);
AND_array_1509 AND_array_1509_c311({a_c[1197:0],311'd0},p_prime[311],c_w_311);
AND_array_1509 AND_array_1509_s311({a_s[1197:0],311'd0},p_prime[311],s_w_311);
AND_array_1509 AND_array_1509_c312({a_c[1196:0],312'd0},p_prime[312],c_w_312);
AND_array_1509 AND_array_1509_s312({a_s[1196:0],312'd0},p_prime[312],s_w_312);
AND_array_1509 AND_array_1509_c313({a_c[1195:0],313'd0},p_prime[313],c_w_313);
AND_array_1509 AND_array_1509_s313({a_s[1195:0],313'd0},p_prime[313],s_w_313);
AND_array_1509 AND_array_1509_c314({a_c[1194:0],314'd0},p_prime[314],c_w_314);
AND_array_1509 AND_array_1509_s314({a_s[1194:0],314'd0},p_prime[314],s_w_314);
AND_array_1509 AND_array_1509_c315({a_c[1193:0],315'd0},p_prime[315],c_w_315);
AND_array_1509 AND_array_1509_s315({a_s[1193:0],315'd0},p_prime[315],s_w_315);
AND_array_1509 AND_array_1509_c316({a_c[1192:0],316'd0},p_prime[316],c_w_316);
AND_array_1509 AND_array_1509_s316({a_s[1192:0],316'd0},p_prime[316],s_w_316);
AND_array_1509 AND_array_1509_c317({a_c[1191:0],317'd0},p_prime[317],c_w_317);
AND_array_1509 AND_array_1509_s317({a_s[1191:0],317'd0},p_prime[317],s_w_317);
AND_array_1509 AND_array_1509_c318({a_c[1190:0],318'd0},p_prime[318],c_w_318);
AND_array_1509 AND_array_1509_s318({a_s[1190:0],318'd0},p_prime[318],s_w_318);
AND_array_1509 AND_array_1509_c319({a_c[1189:0],319'd0},p_prime[319],c_w_319);
AND_array_1509 AND_array_1509_s319({a_s[1189:0],319'd0},p_prime[319],s_w_319);
AND_array_1509 AND_array_1509_c320({a_c[1188:0],320'd0},p_prime[320],c_w_320);
AND_array_1509 AND_array_1509_s320({a_s[1188:0],320'd0},p_prime[320],s_w_320);
AND_array_1509 AND_array_1509_c321({a_c[1187:0],321'd0},p_prime[321],c_w_321);
AND_array_1509 AND_array_1509_s321({a_s[1187:0],321'd0},p_prime[321],s_w_321);
AND_array_1509 AND_array_1509_c322({a_c[1186:0],322'd0},p_prime[322],c_w_322);
AND_array_1509 AND_array_1509_s322({a_s[1186:0],322'd0},p_prime[322],s_w_322);
AND_array_1509 AND_array_1509_c323({a_c[1185:0],323'd0},p_prime[323],c_w_323);
AND_array_1509 AND_array_1509_s323({a_s[1185:0],323'd0},p_prime[323],s_w_323);
AND_array_1509 AND_array_1509_c324({a_c[1184:0],324'd0},p_prime[324],c_w_324);
AND_array_1509 AND_array_1509_s324({a_s[1184:0],324'd0},p_prime[324],s_w_324);
AND_array_1509 AND_array_1509_c325({a_c[1183:0],325'd0},p_prime[325],c_w_325);
AND_array_1509 AND_array_1509_s325({a_s[1183:0],325'd0},p_prime[325],s_w_325);
AND_array_1509 AND_array_1509_c326({a_c[1182:0],326'd0},p_prime[326],c_w_326);
AND_array_1509 AND_array_1509_s326({a_s[1182:0],326'd0},p_prime[326],s_w_326);
AND_array_1509 AND_array_1509_c327({a_c[1181:0],327'd0},p_prime[327],c_w_327);
AND_array_1509 AND_array_1509_s327({a_s[1181:0],327'd0},p_prime[327],s_w_327);
AND_array_1509 AND_array_1509_c328({a_c[1180:0],328'd0},p_prime[328],c_w_328);
AND_array_1509 AND_array_1509_s328({a_s[1180:0],328'd0},p_prime[328],s_w_328);
AND_array_1509 AND_array_1509_c329({a_c[1179:0],329'd0},p_prime[329],c_w_329);
AND_array_1509 AND_array_1509_s329({a_s[1179:0],329'd0},p_prime[329],s_w_329);
AND_array_1509 AND_array_1509_c330({a_c[1178:0],330'd0},p_prime[330],c_w_330);
AND_array_1509 AND_array_1509_s330({a_s[1178:0],330'd0},p_prime[330],s_w_330);
AND_array_1509 AND_array_1509_c331({a_c[1177:0],331'd0},p_prime[331],c_w_331);
AND_array_1509 AND_array_1509_s331({a_s[1177:0],331'd0},p_prime[331],s_w_331);
AND_array_1509 AND_array_1509_c332({a_c[1176:0],332'd0},p_prime[332],c_w_332);
AND_array_1509 AND_array_1509_s332({a_s[1176:0],332'd0},p_prime[332],s_w_332);
AND_array_1509 AND_array_1509_c333({a_c[1175:0],333'd0},p_prime[333],c_w_333);
AND_array_1509 AND_array_1509_s333({a_s[1175:0],333'd0},p_prime[333],s_w_333);
AND_array_1509 AND_array_1509_c334({a_c[1174:0],334'd0},p_prime[334],c_w_334);
AND_array_1509 AND_array_1509_s334({a_s[1174:0],334'd0},p_prime[334],s_w_334);
AND_array_1509 AND_array_1509_c335({a_c[1173:0],335'd0},p_prime[335],c_w_335);
AND_array_1509 AND_array_1509_s335({a_s[1173:0],335'd0},p_prime[335],s_w_335);
AND_array_1509 AND_array_1509_c336({a_c[1172:0],336'd0},p_prime[336],c_w_336);
AND_array_1509 AND_array_1509_s336({a_s[1172:0],336'd0},p_prime[336],s_w_336);
AND_array_1509 AND_array_1509_c337({a_c[1171:0],337'd0},p_prime[337],c_w_337);
AND_array_1509 AND_array_1509_s337({a_s[1171:0],337'd0},p_prime[337],s_w_337);
AND_array_1509 AND_array_1509_c338({a_c[1170:0],338'd0},p_prime[338],c_w_338);
AND_array_1509 AND_array_1509_s338({a_s[1170:0],338'd0},p_prime[338],s_w_338);
AND_array_1509 AND_array_1509_c339({a_c[1169:0],339'd0},p_prime[339],c_w_339);
AND_array_1509 AND_array_1509_s339({a_s[1169:0],339'd0},p_prime[339],s_w_339);
AND_array_1509 AND_array_1509_c340({a_c[1168:0],340'd0},p_prime[340],c_w_340);
AND_array_1509 AND_array_1509_s340({a_s[1168:0],340'd0},p_prime[340],s_w_340);
AND_array_1509 AND_array_1509_c341({a_c[1167:0],341'd0},p_prime[341],c_w_341);
AND_array_1509 AND_array_1509_s341({a_s[1167:0],341'd0},p_prime[341],s_w_341);
AND_array_1509 AND_array_1509_c342({a_c[1166:0],342'd0},p_prime[342],c_w_342);
AND_array_1509 AND_array_1509_s342({a_s[1166:0],342'd0},p_prime[342],s_w_342);
AND_array_1509 AND_array_1509_c343({a_c[1165:0],343'd0},p_prime[343],c_w_343);
AND_array_1509 AND_array_1509_s343({a_s[1165:0],343'd0},p_prime[343],s_w_343);
AND_array_1509 AND_array_1509_c344({a_c[1164:0],344'd0},p_prime[344],c_w_344);
AND_array_1509 AND_array_1509_s344({a_s[1164:0],344'd0},p_prime[344],s_w_344);
AND_array_1509 AND_array_1509_c345({a_c[1163:0],345'd0},p_prime[345],c_w_345);
AND_array_1509 AND_array_1509_s345({a_s[1163:0],345'd0},p_prime[345],s_w_345);
AND_array_1509 AND_array_1509_c346({a_c[1162:0],346'd0},p_prime[346],c_w_346);
AND_array_1509 AND_array_1509_s346({a_s[1162:0],346'd0},p_prime[346],s_w_346);
AND_array_1509 AND_array_1509_c347({a_c[1161:0],347'd0},p_prime[347],c_w_347);
AND_array_1509 AND_array_1509_s347({a_s[1161:0],347'd0},p_prime[347],s_w_347);
AND_array_1509 AND_array_1509_c348({a_c[1160:0],348'd0},p_prime[348],c_w_348);
AND_array_1509 AND_array_1509_s348({a_s[1160:0],348'd0},p_prime[348],s_w_348);
AND_array_1509 AND_array_1509_c349({a_c[1159:0],349'd0},p_prime[349],c_w_349);
AND_array_1509 AND_array_1509_s349({a_s[1159:0],349'd0},p_prime[349],s_w_349);
AND_array_1509 AND_array_1509_c350({a_c[1158:0],350'd0},p_prime[350],c_w_350);
AND_array_1509 AND_array_1509_s350({a_s[1158:0],350'd0},p_prime[350],s_w_350);
AND_array_1509 AND_array_1509_c351({a_c[1157:0],351'd0},p_prime[351],c_w_351);
AND_array_1509 AND_array_1509_s351({a_s[1157:0],351'd0},p_prime[351],s_w_351);
AND_array_1509 AND_array_1509_c352({a_c[1156:0],352'd0},p_prime[352],c_w_352);
AND_array_1509 AND_array_1509_s352({a_s[1156:0],352'd0},p_prime[352],s_w_352);
AND_array_1509 AND_array_1509_c353({a_c[1155:0],353'd0},p_prime[353],c_w_353);
AND_array_1509 AND_array_1509_s353({a_s[1155:0],353'd0},p_prime[353],s_w_353);
AND_array_1509 AND_array_1509_c354({a_c[1154:0],354'd0},p_prime[354],c_w_354);
AND_array_1509 AND_array_1509_s354({a_s[1154:0],354'd0},p_prime[354],s_w_354);
AND_array_1509 AND_array_1509_c355({a_c[1153:0],355'd0},p_prime[355],c_w_355);
AND_array_1509 AND_array_1509_s355({a_s[1153:0],355'd0},p_prime[355],s_w_355);
AND_array_1509 AND_array_1509_c356({a_c[1152:0],356'd0},p_prime[356],c_w_356);
AND_array_1509 AND_array_1509_s356({a_s[1152:0],356'd0},p_prime[356],s_w_356);
AND_array_1509 AND_array_1509_c357({a_c[1151:0],357'd0},p_prime[357],c_w_357);
AND_array_1509 AND_array_1509_s357({a_s[1151:0],357'd0},p_prime[357],s_w_357);
AND_array_1509 AND_array_1509_c358({a_c[1150:0],358'd0},p_prime[358],c_w_358);
AND_array_1509 AND_array_1509_s358({a_s[1150:0],358'd0},p_prime[358],s_w_358);
AND_array_1509 AND_array_1509_c359({a_c[1149:0],359'd0},p_prime[359],c_w_359);
AND_array_1509 AND_array_1509_s359({a_s[1149:0],359'd0},p_prime[359],s_w_359);
AND_array_1509 AND_array_1509_c360({a_c[1148:0],360'd0},p_prime[360],c_w_360);
AND_array_1509 AND_array_1509_s360({a_s[1148:0],360'd0},p_prime[360],s_w_360);
AND_array_1509 AND_array_1509_c361({a_c[1147:0],361'd0},p_prime[361],c_w_361);
AND_array_1509 AND_array_1509_s361({a_s[1147:0],361'd0},p_prime[361],s_w_361);
AND_array_1509 AND_array_1509_c362({a_c[1146:0],362'd0},p_prime[362],c_w_362);
AND_array_1509 AND_array_1509_s362({a_s[1146:0],362'd0},p_prime[362],s_w_362);
AND_array_1509 AND_array_1509_c363({a_c[1145:0],363'd0},p_prime[363],c_w_363);
AND_array_1509 AND_array_1509_s363({a_s[1145:0],363'd0},p_prime[363],s_w_363);
AND_array_1509 AND_array_1509_c364({a_c[1144:0],364'd0},p_prime[364],c_w_364);
AND_array_1509 AND_array_1509_s364({a_s[1144:0],364'd0},p_prime[364],s_w_364);
AND_array_1509 AND_array_1509_c365({a_c[1143:0],365'd0},p_prime[365],c_w_365);
AND_array_1509 AND_array_1509_s365({a_s[1143:0],365'd0},p_prime[365],s_w_365);
AND_array_1509 AND_array_1509_c366({a_c[1142:0],366'd0},p_prime[366],c_w_366);
AND_array_1509 AND_array_1509_s366({a_s[1142:0],366'd0},p_prime[366],s_w_366);
AND_array_1509 AND_array_1509_c367({a_c[1141:0],367'd0},p_prime[367],c_w_367);
AND_array_1509 AND_array_1509_s367({a_s[1141:0],367'd0},p_prime[367],s_w_367);
AND_array_1509 AND_array_1509_c368({a_c[1140:0],368'd0},p_prime[368],c_w_368);
AND_array_1509 AND_array_1509_s368({a_s[1140:0],368'd0},p_prime[368],s_w_368);
AND_array_1509 AND_array_1509_c369({a_c[1139:0],369'd0},p_prime[369],c_w_369);
AND_array_1509 AND_array_1509_s369({a_s[1139:0],369'd0},p_prime[369],s_w_369);
AND_array_1509 AND_array_1509_c370({a_c[1138:0],370'd0},p_prime[370],c_w_370);
AND_array_1509 AND_array_1509_s370({a_s[1138:0],370'd0},p_prime[370],s_w_370);
AND_array_1509 AND_array_1509_c371({a_c[1137:0],371'd0},p_prime[371],c_w_371);
AND_array_1509 AND_array_1509_s371({a_s[1137:0],371'd0},p_prime[371],s_w_371);
AND_array_1509 AND_array_1509_c372({a_c[1136:0],372'd0},p_prime[372],c_w_372);
AND_array_1509 AND_array_1509_s372({a_s[1136:0],372'd0},p_prime[372],s_w_372);
AND_array_1509 AND_array_1509_c373({a_c[1135:0],373'd0},p_prime[373],c_w_373);
AND_array_1509 AND_array_1509_s373({a_s[1135:0],373'd0},p_prime[373],s_w_373);
AND_array_1509 AND_array_1509_c374({a_c[1134:0],374'd0},p_prime[374],c_w_374);
AND_array_1509 AND_array_1509_s374({a_s[1134:0],374'd0},p_prime[374],s_w_374);
AND_array_1509 AND_array_1509_c375({a_c[1133:0],375'd0},p_prime[375],c_w_375);
AND_array_1509 AND_array_1509_s375({a_s[1133:0],375'd0},p_prime[375],s_w_375);
AND_array_1509 AND_array_1509_c376({a_c[1132:0],376'd0},p_prime[376],c_w_376);
AND_array_1509 AND_array_1509_s376({a_s[1132:0],376'd0},p_prime[376],s_w_376);
AND_array_1509 AND_array_1509_c377({a_c[1131:0],377'd0},p_prime[377],c_w_377);
AND_array_1509 AND_array_1509_s377({a_s[1131:0],377'd0},p_prime[377],s_w_377);
AND_array_1509 AND_array_1509_c378({a_c[1130:0],378'd0},p_prime[378],c_w_378);
AND_array_1509 AND_array_1509_s378({a_s[1130:0],378'd0},p_prime[378],s_w_378);
AND_array_1509 AND_array_1509_c379({a_c[1129:0],379'd0},p_prime[379],c_w_379);
AND_array_1509 AND_array_1509_s379({a_s[1129:0],379'd0},p_prime[379],s_w_379);
AND_array_1509 AND_array_1509_c380({a_c[1128:0],380'd0},p_prime[380],c_w_380);
AND_array_1509 AND_array_1509_s380({a_s[1128:0],380'd0},p_prime[380],s_w_380);
AND_array_1509 AND_array_1509_c381({a_c[1127:0],381'd0},p_prime[381],c_w_381);
AND_array_1509 AND_array_1509_s381({a_s[1127:0],381'd0},p_prime[381],s_w_381);
AND_array_1509 AND_array_1509_c382({a_c[1126:0],382'd0},p_prime[382],c_w_382);
AND_array_1509 AND_array_1509_s382({a_s[1126:0],382'd0},p_prime[382],s_w_382);
AND_array_1509 AND_array_1509_c383({a_c[1125:0],383'd0},p_prime[383],c_w_383);
AND_array_1509 AND_array_1509_s383({a_s[1125:0],383'd0},p_prime[383],s_w_383);
AND_array_1509 AND_array_1509_c384({a_c[1124:0],384'd0},p_prime[384],c_w_384);
AND_array_1509 AND_array_1509_s384({a_s[1124:0],384'd0},p_prime[384],s_w_384);
AND_array_1509 AND_array_1509_c385({a_c[1123:0],385'd0},p_prime[385],c_w_385);
AND_array_1509 AND_array_1509_s385({a_s[1123:0],385'd0},p_prime[385],s_w_385);
AND_array_1509 AND_array_1509_c386({a_c[1122:0],386'd0},p_prime[386],c_w_386);
AND_array_1509 AND_array_1509_s386({a_s[1122:0],386'd0},p_prime[386],s_w_386);
AND_array_1509 AND_array_1509_c387({a_c[1121:0],387'd0},p_prime[387],c_w_387);
AND_array_1509 AND_array_1509_s387({a_s[1121:0],387'd0},p_prime[387],s_w_387);
AND_array_1509 AND_array_1509_c388({a_c[1120:0],388'd0},p_prime[388],c_w_388);
AND_array_1509 AND_array_1509_s388({a_s[1120:0],388'd0},p_prime[388],s_w_388);
AND_array_1509 AND_array_1509_c389({a_c[1119:0],389'd0},p_prime[389],c_w_389);
AND_array_1509 AND_array_1509_s389({a_s[1119:0],389'd0},p_prime[389],s_w_389);
AND_array_1509 AND_array_1509_c390({a_c[1118:0],390'd0},p_prime[390],c_w_390);
AND_array_1509 AND_array_1509_s390({a_s[1118:0],390'd0},p_prime[390],s_w_390);
AND_array_1509 AND_array_1509_c391({a_c[1117:0],391'd0},p_prime[391],c_w_391);
AND_array_1509 AND_array_1509_s391({a_s[1117:0],391'd0},p_prime[391],s_w_391);
AND_array_1509 AND_array_1509_c392({a_c[1116:0],392'd0},p_prime[392],c_w_392);
AND_array_1509 AND_array_1509_s392({a_s[1116:0],392'd0},p_prime[392],s_w_392);
AND_array_1509 AND_array_1509_c393({a_c[1115:0],393'd0},p_prime[393],c_w_393);
AND_array_1509 AND_array_1509_s393({a_s[1115:0],393'd0},p_prime[393],s_w_393);
AND_array_1509 AND_array_1509_c394({a_c[1114:0],394'd0},p_prime[394],c_w_394);
AND_array_1509 AND_array_1509_s394({a_s[1114:0],394'd0},p_prime[394],s_w_394);
AND_array_1509 AND_array_1509_c395({a_c[1113:0],395'd0},p_prime[395],c_w_395);
AND_array_1509 AND_array_1509_s395({a_s[1113:0],395'd0},p_prime[395],s_w_395);
AND_array_1509 AND_array_1509_c396({a_c[1112:0],396'd0},p_prime[396],c_w_396);
AND_array_1509 AND_array_1509_s396({a_s[1112:0],396'd0},p_prime[396],s_w_396);
AND_array_1509 AND_array_1509_c397({a_c[1111:0],397'd0},p_prime[397],c_w_397);
AND_array_1509 AND_array_1509_s397({a_s[1111:0],397'd0},p_prime[397],s_w_397);
AND_array_1509 AND_array_1509_c398({a_c[1110:0],398'd0},p_prime[398],c_w_398);
AND_array_1509 AND_array_1509_s398({a_s[1110:0],398'd0},p_prime[398],s_w_398);
AND_array_1509 AND_array_1509_c399({a_c[1109:0],399'd0},p_prime[399],c_w_399);
AND_array_1509 AND_array_1509_s399({a_s[1109:0],399'd0},p_prime[399],s_w_399);
AND_array_1509 AND_array_1509_c400({a_c[1108:0],400'd0},p_prime[400],c_w_400);
AND_array_1509 AND_array_1509_s400({a_s[1108:0],400'd0},p_prime[400],s_w_400);
AND_array_1509 AND_array_1509_c401({a_c[1107:0],401'd0},p_prime[401],c_w_401);
AND_array_1509 AND_array_1509_s401({a_s[1107:0],401'd0},p_prime[401],s_w_401);
AND_array_1509 AND_array_1509_c402({a_c[1106:0],402'd0},p_prime[402],c_w_402);
AND_array_1509 AND_array_1509_s402({a_s[1106:0],402'd0},p_prime[402],s_w_402);
AND_array_1509 AND_array_1509_c403({a_c[1105:0],403'd0},p_prime[403],c_w_403);
AND_array_1509 AND_array_1509_s403({a_s[1105:0],403'd0},p_prime[403],s_w_403);
AND_array_1509 AND_array_1509_c404({a_c[1104:0],404'd0},p_prime[404],c_w_404);
AND_array_1509 AND_array_1509_s404({a_s[1104:0],404'd0},p_prime[404],s_w_404);
AND_array_1509 AND_array_1509_c405({a_c[1103:0],405'd0},p_prime[405],c_w_405);
AND_array_1509 AND_array_1509_s405({a_s[1103:0],405'd0},p_prime[405],s_w_405);
AND_array_1509 AND_array_1509_c406({a_c[1102:0],406'd0},p_prime[406],c_w_406);
AND_array_1509 AND_array_1509_s406({a_s[1102:0],406'd0},p_prime[406],s_w_406);
AND_array_1509 AND_array_1509_c407({a_c[1101:0],407'd0},p_prime[407],c_w_407);
AND_array_1509 AND_array_1509_s407({a_s[1101:0],407'd0},p_prime[407],s_w_407);
AND_array_1509 AND_array_1509_c408({a_c[1100:0],408'd0},p_prime[408],c_w_408);
AND_array_1509 AND_array_1509_s408({a_s[1100:0],408'd0},p_prime[408],s_w_408);
AND_array_1509 AND_array_1509_c409({a_c[1099:0],409'd0},p_prime[409],c_w_409);
AND_array_1509 AND_array_1509_s409({a_s[1099:0],409'd0},p_prime[409],s_w_409);
AND_array_1509 AND_array_1509_c410({a_c[1098:0],410'd0},p_prime[410],c_w_410);
AND_array_1509 AND_array_1509_s410({a_s[1098:0],410'd0},p_prime[410],s_w_410);
AND_array_1509 AND_array_1509_c411({a_c[1097:0],411'd0},p_prime[411],c_w_411);
AND_array_1509 AND_array_1509_s411({a_s[1097:0],411'd0},p_prime[411],s_w_411);
AND_array_1509 AND_array_1509_c412({a_c[1096:0],412'd0},p_prime[412],c_w_412);
AND_array_1509 AND_array_1509_s412({a_s[1096:0],412'd0},p_prime[412],s_w_412);
AND_array_1509 AND_array_1509_c413({a_c[1095:0],413'd0},p_prime[413],c_w_413);
AND_array_1509 AND_array_1509_s413({a_s[1095:0],413'd0},p_prime[413],s_w_413);
AND_array_1509 AND_array_1509_c414({a_c[1094:0],414'd0},p_prime[414],c_w_414);
AND_array_1509 AND_array_1509_s414({a_s[1094:0],414'd0},p_prime[414],s_w_414);
AND_array_1509 AND_array_1509_c415({a_c[1093:0],415'd0},p_prime[415],c_w_415);
AND_array_1509 AND_array_1509_s415({a_s[1093:0],415'd0},p_prime[415],s_w_415);
AND_array_1509 AND_array_1509_c416({a_c[1092:0],416'd0},p_prime[416],c_w_416);
AND_array_1509 AND_array_1509_s416({a_s[1092:0],416'd0},p_prime[416],s_w_416);
AND_array_1509 AND_array_1509_c417({a_c[1091:0],417'd0},p_prime[417],c_w_417);
AND_array_1509 AND_array_1509_s417({a_s[1091:0],417'd0},p_prime[417],s_w_417);
AND_array_1509 AND_array_1509_c418({a_c[1090:0],418'd0},p_prime[418],c_w_418);
AND_array_1509 AND_array_1509_s418({a_s[1090:0],418'd0},p_prime[418],s_w_418);
AND_array_1509 AND_array_1509_c419({a_c[1089:0],419'd0},p_prime[419],c_w_419);
AND_array_1509 AND_array_1509_s419({a_s[1089:0],419'd0},p_prime[419],s_w_419);
AND_array_1509 AND_array_1509_c420({a_c[1088:0],420'd0},p_prime[420],c_w_420);
AND_array_1509 AND_array_1509_s420({a_s[1088:0],420'd0},p_prime[420],s_w_420);
AND_array_1509 AND_array_1509_c421({a_c[1087:0],421'd0},p_prime[421],c_w_421);
AND_array_1509 AND_array_1509_s421({a_s[1087:0],421'd0},p_prime[421],s_w_421);
AND_array_1509 AND_array_1509_c422({a_c[1086:0],422'd0},p_prime[422],c_w_422);
AND_array_1509 AND_array_1509_s422({a_s[1086:0],422'd0},p_prime[422],s_w_422);
AND_array_1509 AND_array_1509_c423({a_c[1085:0],423'd0},p_prime[423],c_w_423);
AND_array_1509 AND_array_1509_s423({a_s[1085:0],423'd0},p_prime[423],s_w_423);
AND_array_1509 AND_array_1509_c424({a_c[1084:0],424'd0},p_prime[424],c_w_424);
AND_array_1509 AND_array_1509_s424({a_s[1084:0],424'd0},p_prime[424],s_w_424);
AND_array_1509 AND_array_1509_c425({a_c[1083:0],425'd0},p_prime[425],c_w_425);
AND_array_1509 AND_array_1509_s425({a_s[1083:0],425'd0},p_prime[425],s_w_425);
AND_array_1509 AND_array_1509_c426({a_c[1082:0],426'd0},p_prime[426],c_w_426);
AND_array_1509 AND_array_1509_s426({a_s[1082:0],426'd0},p_prime[426],s_w_426);
AND_array_1509 AND_array_1509_c427({a_c[1081:0],427'd0},p_prime[427],c_w_427);
AND_array_1509 AND_array_1509_s427({a_s[1081:0],427'd0},p_prime[427],s_w_427);
AND_array_1509 AND_array_1509_c428({a_c[1080:0],428'd0},p_prime[428],c_w_428);
AND_array_1509 AND_array_1509_s428({a_s[1080:0],428'd0},p_prime[428],s_w_428);
AND_array_1509 AND_array_1509_c429({a_c[1079:0],429'd0},p_prime[429],c_w_429);
AND_array_1509 AND_array_1509_s429({a_s[1079:0],429'd0},p_prime[429],s_w_429);
AND_array_1509 AND_array_1509_c430({a_c[1078:0],430'd0},p_prime[430],c_w_430);
AND_array_1509 AND_array_1509_s430({a_s[1078:0],430'd0},p_prime[430],s_w_430);
AND_array_1509 AND_array_1509_c431({a_c[1077:0],431'd0},p_prime[431],c_w_431);
AND_array_1509 AND_array_1509_s431({a_s[1077:0],431'd0},p_prime[431],s_w_431);
AND_array_1509 AND_array_1509_c432({a_c[1076:0],432'd0},p_prime[432],c_w_432);
AND_array_1509 AND_array_1509_s432({a_s[1076:0],432'd0},p_prime[432],s_w_432);
AND_array_1509 AND_array_1509_c433({a_c[1075:0],433'd0},p_prime[433],c_w_433);
AND_array_1509 AND_array_1509_s433({a_s[1075:0],433'd0},p_prime[433],s_w_433);
AND_array_1509 AND_array_1509_c434({a_c[1074:0],434'd0},p_prime[434],c_w_434);
AND_array_1509 AND_array_1509_s434({a_s[1074:0],434'd0},p_prime[434],s_w_434);
AND_array_1509 AND_array_1509_c435({a_c[1073:0],435'd0},p_prime[435],c_w_435);
AND_array_1509 AND_array_1509_s435({a_s[1073:0],435'd0},p_prime[435],s_w_435);
AND_array_1509 AND_array_1509_c436({a_c[1072:0],436'd0},p_prime[436],c_w_436);
AND_array_1509 AND_array_1509_s436({a_s[1072:0],436'd0},p_prime[436],s_w_436);
AND_array_1509 AND_array_1509_c437({a_c[1071:0],437'd0},p_prime[437],c_w_437);
AND_array_1509 AND_array_1509_s437({a_s[1071:0],437'd0},p_prime[437],s_w_437);
AND_array_1509 AND_array_1509_c438({a_c[1070:0],438'd0},p_prime[438],c_w_438);
AND_array_1509 AND_array_1509_s438({a_s[1070:0],438'd0},p_prime[438],s_w_438);
AND_array_1509 AND_array_1509_c439({a_c[1069:0],439'd0},p_prime[439],c_w_439);
AND_array_1509 AND_array_1509_s439({a_s[1069:0],439'd0},p_prime[439],s_w_439);
AND_array_1509 AND_array_1509_c440({a_c[1068:0],440'd0},p_prime[440],c_w_440);
AND_array_1509 AND_array_1509_s440({a_s[1068:0],440'd0},p_prime[440],s_w_440);
AND_array_1509 AND_array_1509_c441({a_c[1067:0],441'd0},p_prime[441],c_w_441);
AND_array_1509 AND_array_1509_s441({a_s[1067:0],441'd0},p_prime[441],s_w_441);
AND_array_1509 AND_array_1509_c442({a_c[1066:0],442'd0},p_prime[442],c_w_442);
AND_array_1509 AND_array_1509_s442({a_s[1066:0],442'd0},p_prime[442],s_w_442);
AND_array_1509 AND_array_1509_c443({a_c[1065:0],443'd0},p_prime[443],c_w_443);
AND_array_1509 AND_array_1509_s443({a_s[1065:0],443'd0},p_prime[443],s_w_443);
AND_array_1509 AND_array_1509_c444({a_c[1064:0],444'd0},p_prime[444],c_w_444);
AND_array_1509 AND_array_1509_s444({a_s[1064:0],444'd0},p_prime[444],s_w_444);
AND_array_1509 AND_array_1509_c445({a_c[1063:0],445'd0},p_prime[445],c_w_445);
AND_array_1509 AND_array_1509_s445({a_s[1063:0],445'd0},p_prime[445],s_w_445);
AND_array_1509 AND_array_1509_c446({a_c[1062:0],446'd0},p_prime[446],c_w_446);
AND_array_1509 AND_array_1509_s446({a_s[1062:0],446'd0},p_prime[446],s_w_446);
AND_array_1509 AND_array_1509_c447({a_c[1061:0],447'd0},p_prime[447],c_w_447);
AND_array_1509 AND_array_1509_s447({a_s[1061:0],447'd0},p_prime[447],s_w_447);
AND_array_1509 AND_array_1509_c448({a_c[1060:0],448'd0},p_prime[448],c_w_448);
AND_array_1509 AND_array_1509_s448({a_s[1060:0],448'd0},p_prime[448],s_w_448);
AND_array_1509 AND_array_1509_c449({a_c[1059:0],449'd0},p_prime[449],c_w_449);
AND_array_1509 AND_array_1509_s449({a_s[1059:0],449'd0},p_prime[449],s_w_449);
AND_array_1509 AND_array_1509_c450({a_c[1058:0],450'd0},p_prime[450],c_w_450);
AND_array_1509 AND_array_1509_s450({a_s[1058:0],450'd0},p_prime[450],s_w_450);
AND_array_1509 AND_array_1509_c451({a_c[1057:0],451'd0},p_prime[451],c_w_451);
AND_array_1509 AND_array_1509_s451({a_s[1057:0],451'd0},p_prime[451],s_w_451);
AND_array_1509 AND_array_1509_c452({a_c[1056:0],452'd0},p_prime[452],c_w_452);
AND_array_1509 AND_array_1509_s452({a_s[1056:0],452'd0},p_prime[452],s_w_452);
AND_array_1509 AND_array_1509_c453({a_c[1055:0],453'd0},p_prime[453],c_w_453);
AND_array_1509 AND_array_1509_s453({a_s[1055:0],453'd0},p_prime[453],s_w_453);
AND_array_1509 AND_array_1509_c454({a_c[1054:0],454'd0},p_prime[454],c_w_454);
AND_array_1509 AND_array_1509_s454({a_s[1054:0],454'd0},p_prime[454],s_w_454);
AND_array_1509 AND_array_1509_c455({a_c[1053:0],455'd0},p_prime[455],c_w_455);
AND_array_1509 AND_array_1509_s455({a_s[1053:0],455'd0},p_prime[455],s_w_455);
AND_array_1509 AND_array_1509_c456({a_c[1052:0],456'd0},p_prime[456],c_w_456);
AND_array_1509 AND_array_1509_s456({a_s[1052:0],456'd0},p_prime[456],s_w_456);
AND_array_1509 AND_array_1509_c457({a_c[1051:0],457'd0},p_prime[457],c_w_457);
AND_array_1509 AND_array_1509_s457({a_s[1051:0],457'd0},p_prime[457],s_w_457);
AND_array_1509 AND_array_1509_c458({a_c[1050:0],458'd0},p_prime[458],c_w_458);
AND_array_1509 AND_array_1509_s458({a_s[1050:0],458'd0},p_prime[458],s_w_458);
AND_array_1509 AND_array_1509_c459({a_c[1049:0],459'd0},p_prime[459],c_w_459);
AND_array_1509 AND_array_1509_s459({a_s[1049:0],459'd0},p_prime[459],s_w_459);
AND_array_1509 AND_array_1509_c460({a_c[1048:0],460'd0},p_prime[460],c_w_460);
AND_array_1509 AND_array_1509_s460({a_s[1048:0],460'd0},p_prime[460],s_w_460);
AND_array_1509 AND_array_1509_c461({a_c[1047:0],461'd0},p_prime[461],c_w_461);
AND_array_1509 AND_array_1509_s461({a_s[1047:0],461'd0},p_prime[461],s_w_461);
AND_array_1509 AND_array_1509_c462({a_c[1046:0],462'd0},p_prime[462],c_w_462);
AND_array_1509 AND_array_1509_s462({a_s[1046:0],462'd0},p_prime[462],s_w_462);
AND_array_1509 AND_array_1509_c463({a_c[1045:0],463'd0},p_prime[463],c_w_463);
AND_array_1509 AND_array_1509_s463({a_s[1045:0],463'd0},p_prime[463],s_w_463);
AND_array_1509 AND_array_1509_c464({a_c[1044:0],464'd0},p_prime[464],c_w_464);
AND_array_1509 AND_array_1509_s464({a_s[1044:0],464'd0},p_prime[464],s_w_464);
AND_array_1509 AND_array_1509_c465({a_c[1043:0],465'd0},p_prime[465],c_w_465);
AND_array_1509 AND_array_1509_s465({a_s[1043:0],465'd0},p_prime[465],s_w_465);
AND_array_1509 AND_array_1509_c466({a_c[1042:0],466'd0},p_prime[466],c_w_466);
AND_array_1509 AND_array_1509_s466({a_s[1042:0],466'd0},p_prime[466],s_w_466);
AND_array_1509 AND_array_1509_c467({a_c[1041:0],467'd0},p_prime[467],c_w_467);
AND_array_1509 AND_array_1509_s467({a_s[1041:0],467'd0},p_prime[467],s_w_467);
AND_array_1509 AND_array_1509_c468({a_c[1040:0],468'd0},p_prime[468],c_w_468);
AND_array_1509 AND_array_1509_s468({a_s[1040:0],468'd0},p_prime[468],s_w_468);
AND_array_1509 AND_array_1509_c469({a_c[1039:0],469'd0},p_prime[469],c_w_469);
AND_array_1509 AND_array_1509_s469({a_s[1039:0],469'd0},p_prime[469],s_w_469);
AND_array_1509 AND_array_1509_c470({a_c[1038:0],470'd0},p_prime[470],c_w_470);
AND_array_1509 AND_array_1509_s470({a_s[1038:0],470'd0},p_prime[470],s_w_470);
AND_array_1509 AND_array_1509_c471({a_c[1037:0],471'd0},p_prime[471],c_w_471);
AND_array_1509 AND_array_1509_s471({a_s[1037:0],471'd0},p_prime[471],s_w_471);
AND_array_1509 AND_array_1509_c472({a_c[1036:0],472'd0},p_prime[472],c_w_472);
AND_array_1509 AND_array_1509_s472({a_s[1036:0],472'd0},p_prime[472],s_w_472);
AND_array_1509 AND_array_1509_c473({a_c[1035:0],473'd0},p_prime[473],c_w_473);
AND_array_1509 AND_array_1509_s473({a_s[1035:0],473'd0},p_prime[473],s_w_473);
AND_array_1509 AND_array_1509_c474({a_c[1034:0],474'd0},p_prime[474],c_w_474);
AND_array_1509 AND_array_1509_s474({a_s[1034:0],474'd0},p_prime[474],s_w_474);
AND_array_1509 AND_array_1509_c475({a_c[1033:0],475'd0},p_prime[475],c_w_475);
AND_array_1509 AND_array_1509_s475({a_s[1033:0],475'd0},p_prime[475],s_w_475);
AND_array_1509 AND_array_1509_c476({a_c[1032:0],476'd0},p_prime[476],c_w_476);
AND_array_1509 AND_array_1509_s476({a_s[1032:0],476'd0},p_prime[476],s_w_476);
AND_array_1509 AND_array_1509_c477({a_c[1031:0],477'd0},p_prime[477],c_w_477);
AND_array_1509 AND_array_1509_s477({a_s[1031:0],477'd0},p_prime[477],s_w_477);
AND_array_1509 AND_array_1509_c478({a_c[1030:0],478'd0},p_prime[478],c_w_478);
AND_array_1509 AND_array_1509_s478({a_s[1030:0],478'd0},p_prime[478],s_w_478);
AND_array_1509 AND_array_1509_c479({a_c[1029:0],479'd0},p_prime[479],c_w_479);
AND_array_1509 AND_array_1509_s479({a_s[1029:0],479'd0},p_prime[479],s_w_479);
AND_array_1509 AND_array_1509_c480({a_c[1028:0],480'd0},p_prime[480],c_w_480);
AND_array_1509 AND_array_1509_s480({a_s[1028:0],480'd0},p_prime[480],s_w_480);
AND_array_1509 AND_array_1509_c481({a_c[1027:0],481'd0},p_prime[481],c_w_481);
AND_array_1509 AND_array_1509_s481({a_s[1027:0],481'd0},p_prime[481],s_w_481);
AND_array_1509 AND_array_1509_c482({a_c[1026:0],482'd0},p_prime[482],c_w_482);
AND_array_1509 AND_array_1509_s482({a_s[1026:0],482'd0},p_prime[482],s_w_482);
AND_array_1509 AND_array_1509_c483({a_c[1025:0],483'd0},p_prime[483],c_w_483);
AND_array_1509 AND_array_1509_s483({a_s[1025:0],483'd0},p_prime[483],s_w_483);
AND_array_1509 AND_array_1509_c484({a_c[1024:0],484'd0},p_prime[484],c_w_484);
AND_array_1509 AND_array_1509_s484({a_s[1024:0],484'd0},p_prime[484],s_w_484);
AND_array_1509 AND_array_1509_c485({a_c[1023:0],485'd0},p_prime[485],c_w_485);
AND_array_1509 AND_array_1509_s485({a_s[1023:0],485'd0},p_prime[485],s_w_485);
AND_array_1509 AND_array_1509_c486({a_c[1022:0],486'd0},p_prime[486],c_w_486);
AND_array_1509 AND_array_1509_s486({a_s[1022:0],486'd0},p_prime[486],s_w_486);
AND_array_1509 AND_array_1509_c487({a_c[1021:0],487'd0},p_prime[487],c_w_487);
AND_array_1509 AND_array_1509_s487({a_s[1021:0],487'd0},p_prime[487],s_w_487);
AND_array_1509 AND_array_1509_c488({a_c[1020:0],488'd0},p_prime[488],c_w_488);
AND_array_1509 AND_array_1509_s488({a_s[1020:0],488'd0},p_prime[488],s_w_488);
AND_array_1509 AND_array_1509_c489({a_c[1019:0],489'd0},p_prime[489],c_w_489);
AND_array_1509 AND_array_1509_s489({a_s[1019:0],489'd0},p_prime[489],s_w_489);
AND_array_1509 AND_array_1509_c490({a_c[1018:0],490'd0},p_prime[490],c_w_490);
AND_array_1509 AND_array_1509_s490({a_s[1018:0],490'd0},p_prime[490],s_w_490);
AND_array_1509 AND_array_1509_c491({a_c[1017:0],491'd0},p_prime[491],c_w_491);
AND_array_1509 AND_array_1509_s491({a_s[1017:0],491'd0},p_prime[491],s_w_491);
AND_array_1509 AND_array_1509_c492({a_c[1016:0],492'd0},p_prime[492],c_w_492);
AND_array_1509 AND_array_1509_s492({a_s[1016:0],492'd0},p_prime[492],s_w_492);
AND_array_1509 AND_array_1509_c493({a_c[1015:0],493'd0},p_prime[493],c_w_493);
AND_array_1509 AND_array_1509_s493({a_s[1015:0],493'd0},p_prime[493],s_w_493);
AND_array_1509 AND_array_1509_c494({a_c[1014:0],494'd0},p_prime[494],c_w_494);
AND_array_1509 AND_array_1509_s494({a_s[1014:0],494'd0},p_prime[494],s_w_494);
AND_array_1509 AND_array_1509_c495({a_c[1013:0],495'd0},p_prime[495],c_w_495);
AND_array_1509 AND_array_1509_s495({a_s[1013:0],495'd0},p_prime[495],s_w_495);
AND_array_1509 AND_array_1509_c496({a_c[1012:0],496'd0},p_prime[496],c_w_496);
AND_array_1509 AND_array_1509_s496({a_s[1012:0],496'd0},p_prime[496],s_w_496);
AND_array_1509 AND_array_1509_c497({a_c[1011:0],497'd0},p_prime[497],c_w_497);
AND_array_1509 AND_array_1509_s497({a_s[1011:0],497'd0},p_prime[497],s_w_497);
AND_array_1509 AND_array_1509_c498({a_c[1010:0],498'd0},p_prime[498],c_w_498);
AND_array_1509 AND_array_1509_s498({a_s[1010:0],498'd0},p_prime[498],s_w_498);
AND_array_1509 AND_array_1509_c499({a_c[1009:0],499'd0},p_prime[499],c_w_499);
AND_array_1509 AND_array_1509_s499({a_s[1009:0],499'd0},p_prime[499],s_w_499);
AND_array_1509 AND_array_1509_c500({a_c[1008:0],500'd0},p_prime[500],c_w_500);
AND_array_1509 AND_array_1509_s500({a_s[1008:0],500'd0},p_prime[500],s_w_500);
AND_array_1509 AND_array_1509_c501({a_c[1007:0],501'd0},p_prime[501],c_w_501);
AND_array_1509 AND_array_1509_s501({a_s[1007:0],501'd0},p_prime[501],s_w_501);
AND_array_1509 AND_array_1509_c502({a_c[1006:0],502'd0},p_prime[502],c_w_502);
AND_array_1509 AND_array_1509_s502({a_s[1006:0],502'd0},p_prime[502],s_w_502);
AND_array_1509 AND_array_1509_c503({a_c[1005:0],503'd0},p_prime[503],c_w_503);
AND_array_1509 AND_array_1509_s503({a_s[1005:0],503'd0},p_prime[503],s_w_503);
AND_array_1509 AND_array_1509_c504({a_c[1004:0],504'd0},p_prime[504],c_w_504);
AND_array_1509 AND_array_1509_s504({a_s[1004:0],504'd0},p_prime[504],s_w_504);
AND_array_1509 AND_array_1509_c505({a_c[1003:0],505'd0},p_prime[505],c_w_505);
AND_array_1509 AND_array_1509_s505({a_s[1003:0],505'd0},p_prime[505],s_w_505);
AND_array_1509 AND_array_1509_c506({a_c[1002:0],506'd0},p_prime[506],c_w_506);
AND_array_1509 AND_array_1509_s506({a_s[1002:0],506'd0},p_prime[506],s_w_506);
AND_array_1509 AND_array_1509_c507({a_c[1001:0],507'd0},p_prime[507],c_w_507);
AND_array_1509 AND_array_1509_s507({a_s[1001:0],507'd0},p_prime[507],s_w_507);
AND_array_1509 AND_array_1509_c508({a_c[1000:0],508'd0},p_prime[508],c_w_508);
AND_array_1509 AND_array_1509_s508({a_s[1000:0],508'd0},p_prime[508],s_w_508);
AND_array_1509 AND_array_1509_c509({a_c[999:0],509'd0},p_prime[509],c_w_509);
AND_array_1509 AND_array_1509_s509({a_s[999:0],509'd0},p_prime[509],s_w_509);
AND_array_1509 AND_array_1509_c510({a_c[998:0],510'd0},p_prime[510],c_w_510);
AND_array_1509 AND_array_1509_s510({a_s[998:0],510'd0},p_prime[510],s_w_510);
AND_array_1509 AND_array_1509_c511({a_c[997:0],511'd0},p_prime[511],c_w_511);
AND_array_1509 AND_array_1509_s511({a_s[997:0],511'd0},p_prime[511],s_w_511);
AND_array_1509 AND_array_1509_c512({a_c[996:0],512'd0},p_prime[512],c_w_512);
AND_array_1509 AND_array_1509_s512({a_s[996:0],512'd0},p_prime[512],s_w_512);
AND_array_1509 AND_array_1509_c513({a_c[995:0],513'd0},p_prime[513],c_w_513);
AND_array_1509 AND_array_1509_s513({a_s[995:0],513'd0},p_prime[513],s_w_513);
AND_array_1509 AND_array_1509_c514({a_c[994:0],514'd0},p_prime[514],c_w_514);
AND_array_1509 AND_array_1509_s514({a_s[994:0],514'd0},p_prime[514],s_w_514);
AND_array_1509 AND_array_1509_c515({a_c[993:0],515'd0},p_prime[515],c_w_515);
AND_array_1509 AND_array_1509_s515({a_s[993:0],515'd0},p_prime[515],s_w_515);
AND_array_1509 AND_array_1509_c516({a_c[992:0],516'd0},p_prime[516],c_w_516);
AND_array_1509 AND_array_1509_s516({a_s[992:0],516'd0},p_prime[516],s_w_516);
AND_array_1509 AND_array_1509_c517({a_c[991:0],517'd0},p_prime[517],c_w_517);
AND_array_1509 AND_array_1509_s517({a_s[991:0],517'd0},p_prime[517],s_w_517);
AND_array_1509 AND_array_1509_c518({a_c[990:0],518'd0},p_prime[518],c_w_518);
AND_array_1509 AND_array_1509_s518({a_s[990:0],518'd0},p_prime[518],s_w_518);
AND_array_1509 AND_array_1509_c519({a_c[989:0],519'd0},p_prime[519],c_w_519);
AND_array_1509 AND_array_1509_s519({a_s[989:0],519'd0},p_prime[519],s_w_519);
AND_array_1509 AND_array_1509_c520({a_c[988:0],520'd0},p_prime[520],c_w_520);
AND_array_1509 AND_array_1509_s520({a_s[988:0],520'd0},p_prime[520],s_w_520);
AND_array_1509 AND_array_1509_c521({a_c[987:0],521'd0},p_prime[521],c_w_521);
AND_array_1509 AND_array_1509_s521({a_s[987:0],521'd0},p_prime[521],s_w_521);
AND_array_1509 AND_array_1509_c522({a_c[986:0],522'd0},p_prime[522],c_w_522);
AND_array_1509 AND_array_1509_s522({a_s[986:0],522'd0},p_prime[522],s_w_522);
AND_array_1509 AND_array_1509_c523({a_c[985:0],523'd0},p_prime[523],c_w_523);
AND_array_1509 AND_array_1509_s523({a_s[985:0],523'd0},p_prime[523],s_w_523);
AND_array_1509 AND_array_1509_c524({a_c[984:0],524'd0},p_prime[524],c_w_524);
AND_array_1509 AND_array_1509_s524({a_s[984:0],524'd0},p_prime[524],s_w_524);
AND_array_1509 AND_array_1509_c525({a_c[983:0],525'd0},p_prime[525],c_w_525);
AND_array_1509 AND_array_1509_s525({a_s[983:0],525'd0},p_prime[525],s_w_525);
AND_array_1509 AND_array_1509_c526({a_c[982:0],526'd0},p_prime[526],c_w_526);
AND_array_1509 AND_array_1509_s526({a_s[982:0],526'd0},p_prime[526],s_w_526);
AND_array_1509 AND_array_1509_c527({a_c[981:0],527'd0},p_prime[527],c_w_527);
AND_array_1509 AND_array_1509_s527({a_s[981:0],527'd0},p_prime[527],s_w_527);
AND_array_1509 AND_array_1509_c528({a_c[980:0],528'd0},p_prime[528],c_w_528);
AND_array_1509 AND_array_1509_s528({a_s[980:0],528'd0},p_prime[528],s_w_528);
AND_array_1509 AND_array_1509_c529({a_c[979:0],529'd0},p_prime[529],c_w_529);
AND_array_1509 AND_array_1509_s529({a_s[979:0],529'd0},p_prime[529],s_w_529);
AND_array_1509 AND_array_1509_c530({a_c[978:0],530'd0},p_prime[530],c_w_530);
AND_array_1509 AND_array_1509_s530({a_s[978:0],530'd0},p_prime[530],s_w_530);
AND_array_1509 AND_array_1509_c531({a_c[977:0],531'd0},p_prime[531],c_w_531);
AND_array_1509 AND_array_1509_s531({a_s[977:0],531'd0},p_prime[531],s_w_531);
AND_array_1509 AND_array_1509_c532({a_c[976:0],532'd0},p_prime[532],c_w_532);
AND_array_1509 AND_array_1509_s532({a_s[976:0],532'd0},p_prime[532],s_w_532);
AND_array_1509 AND_array_1509_c533({a_c[975:0],533'd0},p_prime[533],c_w_533);
AND_array_1509 AND_array_1509_s533({a_s[975:0],533'd0},p_prime[533],s_w_533);
AND_array_1509 AND_array_1509_c534({a_c[974:0],534'd0},p_prime[534],c_w_534);
AND_array_1509 AND_array_1509_s534({a_s[974:0],534'd0},p_prime[534],s_w_534);
AND_array_1509 AND_array_1509_c535({a_c[973:0],535'd0},p_prime[535],c_w_535);
AND_array_1509 AND_array_1509_s535({a_s[973:0],535'd0},p_prime[535],s_w_535);
AND_array_1509 AND_array_1509_c536({a_c[972:0],536'd0},p_prime[536],c_w_536);
AND_array_1509 AND_array_1509_s536({a_s[972:0],536'd0},p_prime[536],s_w_536);
AND_array_1509 AND_array_1509_c537({a_c[971:0],537'd0},p_prime[537],c_w_537);
AND_array_1509 AND_array_1509_s537({a_s[971:0],537'd0},p_prime[537],s_w_537);
AND_array_1509 AND_array_1509_c538({a_c[970:0],538'd0},p_prime[538],c_w_538);
AND_array_1509 AND_array_1509_s538({a_s[970:0],538'd0},p_prime[538],s_w_538);
AND_array_1509 AND_array_1509_c539({a_c[969:0],539'd0},p_prime[539],c_w_539);
AND_array_1509 AND_array_1509_s539({a_s[969:0],539'd0},p_prime[539],s_w_539);
AND_array_1509 AND_array_1509_c540({a_c[968:0],540'd0},p_prime[540],c_w_540);
AND_array_1509 AND_array_1509_s540({a_s[968:0],540'd0},p_prime[540],s_w_540);
AND_array_1509 AND_array_1509_c541({a_c[967:0],541'd0},p_prime[541],c_w_541);
AND_array_1509 AND_array_1509_s541({a_s[967:0],541'd0},p_prime[541],s_w_541);
AND_array_1509 AND_array_1509_c542({a_c[966:0],542'd0},p_prime[542],c_w_542);
AND_array_1509 AND_array_1509_s542({a_s[966:0],542'd0},p_prime[542],s_w_542);
AND_array_1509 AND_array_1509_c543({a_c[965:0],543'd0},p_prime[543],c_w_543);
AND_array_1509 AND_array_1509_s543({a_s[965:0],543'd0},p_prime[543],s_w_543);
AND_array_1509 AND_array_1509_c544({a_c[964:0],544'd0},p_prime[544],c_w_544);
AND_array_1509 AND_array_1509_s544({a_s[964:0],544'd0},p_prime[544],s_w_544);
AND_array_1509 AND_array_1509_c545({a_c[963:0],545'd0},p_prime[545],c_w_545);
AND_array_1509 AND_array_1509_s545({a_s[963:0],545'd0},p_prime[545],s_w_545);
AND_array_1509 AND_array_1509_c546({a_c[962:0],546'd0},p_prime[546],c_w_546);
AND_array_1509 AND_array_1509_s546({a_s[962:0],546'd0},p_prime[546],s_w_546);
AND_array_1509 AND_array_1509_c547({a_c[961:0],547'd0},p_prime[547],c_w_547);
AND_array_1509 AND_array_1509_s547({a_s[961:0],547'd0},p_prime[547],s_w_547);
AND_array_1509 AND_array_1509_c548({a_c[960:0],548'd0},p_prime[548],c_w_548);
AND_array_1509 AND_array_1509_s548({a_s[960:0],548'd0},p_prime[548],s_w_548);
AND_array_1509 AND_array_1509_c549({a_c[959:0],549'd0},p_prime[549],c_w_549);
AND_array_1509 AND_array_1509_s549({a_s[959:0],549'd0},p_prime[549],s_w_549);
AND_array_1509 AND_array_1509_c550({a_c[958:0],550'd0},p_prime[550],c_w_550);
AND_array_1509 AND_array_1509_s550({a_s[958:0],550'd0},p_prime[550],s_w_550);
AND_array_1509 AND_array_1509_c551({a_c[957:0],551'd0},p_prime[551],c_w_551);
AND_array_1509 AND_array_1509_s551({a_s[957:0],551'd0},p_prime[551],s_w_551);
AND_array_1509 AND_array_1509_c552({a_c[956:0],552'd0},p_prime[552],c_w_552);
AND_array_1509 AND_array_1509_s552({a_s[956:0],552'd0},p_prime[552],s_w_552);
AND_array_1509 AND_array_1509_c553({a_c[955:0],553'd0},p_prime[553],c_w_553);
AND_array_1509 AND_array_1509_s553({a_s[955:0],553'd0},p_prime[553],s_w_553);
AND_array_1509 AND_array_1509_c554({a_c[954:0],554'd0},p_prime[554],c_w_554);
AND_array_1509 AND_array_1509_s554({a_s[954:0],554'd0},p_prime[554],s_w_554);
AND_array_1509 AND_array_1509_c555({a_c[953:0],555'd0},p_prime[555],c_w_555);
AND_array_1509 AND_array_1509_s555({a_s[953:0],555'd0},p_prime[555],s_w_555);
AND_array_1509 AND_array_1509_c556({a_c[952:0],556'd0},p_prime[556],c_w_556);
AND_array_1509 AND_array_1509_s556({a_s[952:0],556'd0},p_prime[556],s_w_556);
AND_array_1509 AND_array_1509_c557({a_c[951:0],557'd0},p_prime[557],c_w_557);
AND_array_1509 AND_array_1509_s557({a_s[951:0],557'd0},p_prime[557],s_w_557);
AND_array_1509 AND_array_1509_c558({a_c[950:0],558'd0},p_prime[558],c_w_558);
AND_array_1509 AND_array_1509_s558({a_s[950:0],558'd0},p_prime[558],s_w_558);
AND_array_1509 AND_array_1509_c559({a_c[949:0],559'd0},p_prime[559],c_w_559);
AND_array_1509 AND_array_1509_s559({a_s[949:0],559'd0},p_prime[559],s_w_559);
AND_array_1509 AND_array_1509_c560({a_c[948:0],560'd0},p_prime[560],c_w_560);
AND_array_1509 AND_array_1509_s560({a_s[948:0],560'd0},p_prime[560],s_w_560);
AND_array_1509 AND_array_1509_c561({a_c[947:0],561'd0},p_prime[561],c_w_561);
AND_array_1509 AND_array_1509_s561({a_s[947:0],561'd0},p_prime[561],s_w_561);
AND_array_1509 AND_array_1509_c562({a_c[946:0],562'd0},p_prime[562],c_w_562);
AND_array_1509 AND_array_1509_s562({a_s[946:0],562'd0},p_prime[562],s_w_562);
AND_array_1509 AND_array_1509_c563({a_c[945:0],563'd0},p_prime[563],c_w_563);
AND_array_1509 AND_array_1509_s563({a_s[945:0],563'd0},p_prime[563],s_w_563);
AND_array_1509 AND_array_1509_c564({a_c[944:0],564'd0},p_prime[564],c_w_564);
AND_array_1509 AND_array_1509_s564({a_s[944:0],564'd0},p_prime[564],s_w_564);
AND_array_1509 AND_array_1509_c565({a_c[943:0],565'd0},p_prime[565],c_w_565);
AND_array_1509 AND_array_1509_s565({a_s[943:0],565'd0},p_prime[565],s_w_565);
AND_array_1509 AND_array_1509_c566({a_c[942:0],566'd0},p_prime[566],c_w_566);
AND_array_1509 AND_array_1509_s566({a_s[942:0],566'd0},p_prime[566],s_w_566);
AND_array_1509 AND_array_1509_c567({a_c[941:0],567'd0},p_prime[567],c_w_567);
AND_array_1509 AND_array_1509_s567({a_s[941:0],567'd0},p_prime[567],s_w_567);
AND_array_1509 AND_array_1509_c568({a_c[940:0],568'd0},p_prime[568],c_w_568);
AND_array_1509 AND_array_1509_s568({a_s[940:0],568'd0},p_prime[568],s_w_568);
AND_array_1509 AND_array_1509_c569({a_c[939:0],569'd0},p_prime[569],c_w_569);
AND_array_1509 AND_array_1509_s569({a_s[939:0],569'd0},p_prime[569],s_w_569);
AND_array_1509 AND_array_1509_c570({a_c[938:0],570'd0},p_prime[570],c_w_570);
AND_array_1509 AND_array_1509_s570({a_s[938:0],570'd0},p_prime[570],s_w_570);
AND_array_1509 AND_array_1509_c571({a_c[937:0],571'd0},p_prime[571],c_w_571);
AND_array_1509 AND_array_1509_s571({a_s[937:0],571'd0},p_prime[571],s_w_571);
AND_array_1509 AND_array_1509_c572({a_c[936:0],572'd0},p_prime[572],c_w_572);
AND_array_1509 AND_array_1509_s572({a_s[936:0],572'd0},p_prime[572],s_w_572);
AND_array_1509 AND_array_1509_c573({a_c[935:0],573'd0},p_prime[573],c_w_573);
AND_array_1509 AND_array_1509_s573({a_s[935:0],573'd0},p_prime[573],s_w_573);
AND_array_1509 AND_array_1509_c574({a_c[934:0],574'd0},p_prime[574],c_w_574);
AND_array_1509 AND_array_1509_s574({a_s[934:0],574'd0},p_prime[574],s_w_574);
AND_array_1509 AND_array_1509_c575({a_c[933:0],575'd0},p_prime[575],c_w_575);
AND_array_1509 AND_array_1509_s575({a_s[933:0],575'd0},p_prime[575],s_w_575);
AND_array_1509 AND_array_1509_c576({a_c[932:0],576'd0},p_prime[576],c_w_576);
AND_array_1509 AND_array_1509_s576({a_s[932:0],576'd0},p_prime[576],s_w_576);
AND_array_1509 AND_array_1509_c577({a_c[931:0],577'd0},p_prime[577],c_w_577);
AND_array_1509 AND_array_1509_s577({a_s[931:0],577'd0},p_prime[577],s_w_577);
AND_array_1509 AND_array_1509_c578({a_c[930:0],578'd0},p_prime[578],c_w_578);
AND_array_1509 AND_array_1509_s578({a_s[930:0],578'd0},p_prime[578],s_w_578);
AND_array_1509 AND_array_1509_c579({a_c[929:0],579'd0},p_prime[579],c_w_579);
AND_array_1509 AND_array_1509_s579({a_s[929:0],579'd0},p_prime[579],s_w_579);
AND_array_1509 AND_array_1509_c580({a_c[928:0],580'd0},p_prime[580],c_w_580);
AND_array_1509 AND_array_1509_s580({a_s[928:0],580'd0},p_prime[580],s_w_580);
AND_array_1509 AND_array_1509_c581({a_c[927:0],581'd0},p_prime[581],c_w_581);
AND_array_1509 AND_array_1509_s581({a_s[927:0],581'd0},p_prime[581],s_w_581);
AND_array_1509 AND_array_1509_c582({a_c[926:0],582'd0},p_prime[582],c_w_582);
AND_array_1509 AND_array_1509_s582({a_s[926:0],582'd0},p_prime[582],s_w_582);
AND_array_1509 AND_array_1509_c583({a_c[925:0],583'd0},p_prime[583],c_w_583);
AND_array_1509 AND_array_1509_s583({a_s[925:0],583'd0},p_prime[583],s_w_583);
AND_array_1509 AND_array_1509_c584({a_c[924:0],584'd0},p_prime[584],c_w_584);
AND_array_1509 AND_array_1509_s584({a_s[924:0],584'd0},p_prime[584],s_w_584);
AND_array_1509 AND_array_1509_c585({a_c[923:0],585'd0},p_prime[585],c_w_585);
AND_array_1509 AND_array_1509_s585({a_s[923:0],585'd0},p_prime[585],s_w_585);
AND_array_1509 AND_array_1509_c586({a_c[922:0],586'd0},p_prime[586],c_w_586);
AND_array_1509 AND_array_1509_s586({a_s[922:0],586'd0},p_prime[586],s_w_586);
AND_array_1509 AND_array_1509_c587({a_c[921:0],587'd0},p_prime[587],c_w_587);
AND_array_1509 AND_array_1509_s587({a_s[921:0],587'd0},p_prime[587],s_w_587);
AND_array_1509 AND_array_1509_c588({a_c[920:0],588'd0},p_prime[588],c_w_588);
AND_array_1509 AND_array_1509_s588({a_s[920:0],588'd0},p_prime[588],s_w_588);
AND_array_1509 AND_array_1509_c589({a_c[919:0],589'd0},p_prime[589],c_w_589);
AND_array_1509 AND_array_1509_s589({a_s[919:0],589'd0},p_prime[589],s_w_589);
AND_array_1509 AND_array_1509_c590({a_c[918:0],590'd0},p_prime[590],c_w_590);
AND_array_1509 AND_array_1509_s590({a_s[918:0],590'd0},p_prime[590],s_w_590);
AND_array_1509 AND_array_1509_c591({a_c[917:0],591'd0},p_prime[591],c_w_591);
AND_array_1509 AND_array_1509_s591({a_s[917:0],591'd0},p_prime[591],s_w_591);
AND_array_1509 AND_array_1509_c592({a_c[916:0],592'd0},p_prime[592],c_w_592);
AND_array_1509 AND_array_1509_s592({a_s[916:0],592'd0},p_prime[592],s_w_592);
AND_array_1509 AND_array_1509_c593({a_c[915:0],593'd0},p_prime[593],c_w_593);
AND_array_1509 AND_array_1509_s593({a_s[915:0],593'd0},p_prime[593],s_w_593);
AND_array_1509 AND_array_1509_c594({a_c[914:0],594'd0},p_prime[594],c_w_594);
AND_array_1509 AND_array_1509_s594({a_s[914:0],594'd0},p_prime[594],s_w_594);
AND_array_1509 AND_array_1509_c595({a_c[913:0],595'd0},p_prime[595],c_w_595);
AND_array_1509 AND_array_1509_s595({a_s[913:0],595'd0},p_prime[595],s_w_595);
AND_array_1509 AND_array_1509_c596({a_c[912:0],596'd0},p_prime[596],c_w_596);
AND_array_1509 AND_array_1509_s596({a_s[912:0],596'd0},p_prime[596],s_w_596);
AND_array_1509 AND_array_1509_c597({a_c[911:0],597'd0},p_prime[597],c_w_597);
AND_array_1509 AND_array_1509_s597({a_s[911:0],597'd0},p_prime[597],s_w_597);
AND_array_1509 AND_array_1509_c598({a_c[910:0],598'd0},p_prime[598],c_w_598);
AND_array_1509 AND_array_1509_s598({a_s[910:0],598'd0},p_prime[598],s_w_598);
AND_array_1509 AND_array_1509_c599({a_c[909:0],599'd0},p_prime[599],c_w_599);
AND_array_1509 AND_array_1509_s599({a_s[909:0],599'd0},p_prime[599],s_w_599);
AND_array_1509 AND_array_1509_c600({a_c[908:0],600'd0},p_prime[600],c_w_600);
AND_array_1509 AND_array_1509_s600({a_s[908:0],600'd0},p_prime[600],s_w_600);
AND_array_1509 AND_array_1509_c601({a_c[907:0],601'd0},p_prime[601],c_w_601);
AND_array_1509 AND_array_1509_s601({a_s[907:0],601'd0},p_prime[601],s_w_601);
AND_array_1509 AND_array_1509_c602({a_c[906:0],602'd0},p_prime[602],c_w_602);
AND_array_1509 AND_array_1509_s602({a_s[906:0],602'd0},p_prime[602],s_w_602);
AND_array_1509 AND_array_1509_c603({a_c[905:0],603'd0},p_prime[603],c_w_603);
AND_array_1509 AND_array_1509_s603({a_s[905:0],603'd0},p_prime[603],s_w_603);
AND_array_1509 AND_array_1509_c604({a_c[904:0],604'd0},p_prime[604],c_w_604);
AND_array_1509 AND_array_1509_s604({a_s[904:0],604'd0},p_prime[604],s_w_604);
AND_array_1509 AND_array_1509_c605({a_c[903:0],605'd0},p_prime[605],c_w_605);
AND_array_1509 AND_array_1509_s605({a_s[903:0],605'd0},p_prime[605],s_w_605);
AND_array_1509 AND_array_1509_c606({a_c[902:0],606'd0},p_prime[606],c_w_606);
AND_array_1509 AND_array_1509_s606({a_s[902:0],606'd0},p_prime[606],s_w_606);
AND_array_1509 AND_array_1509_c607({a_c[901:0],607'd0},p_prime[607],c_w_607);
AND_array_1509 AND_array_1509_s607({a_s[901:0],607'd0},p_prime[607],s_w_607);
AND_array_1509 AND_array_1509_c608({a_c[900:0],608'd0},p_prime[608],c_w_608);
AND_array_1509 AND_array_1509_s608({a_s[900:0],608'd0},p_prime[608],s_w_608);
AND_array_1509 AND_array_1509_c609({a_c[899:0],609'd0},p_prime[609],c_w_609);
AND_array_1509 AND_array_1509_s609({a_s[899:0],609'd0},p_prime[609],s_w_609);
AND_array_1509 AND_array_1509_c610({a_c[898:0],610'd0},p_prime[610],c_w_610);
AND_array_1509 AND_array_1509_s610({a_s[898:0],610'd0},p_prime[610],s_w_610);
AND_array_1509 AND_array_1509_c611({a_c[897:0],611'd0},p_prime[611],c_w_611);
AND_array_1509 AND_array_1509_s611({a_s[897:0],611'd0},p_prime[611],s_w_611);
AND_array_1509 AND_array_1509_c612({a_c[896:0],612'd0},p_prime[612],c_w_612);
AND_array_1509 AND_array_1509_s612({a_s[896:0],612'd0},p_prime[612],s_w_612);
AND_array_1509 AND_array_1509_c613({a_c[895:0],613'd0},p_prime[613],c_w_613);
AND_array_1509 AND_array_1509_s613({a_s[895:0],613'd0},p_prime[613],s_w_613);
AND_array_1509 AND_array_1509_c614({a_c[894:0],614'd0},p_prime[614],c_w_614);
AND_array_1509 AND_array_1509_s614({a_s[894:0],614'd0},p_prime[614],s_w_614);
AND_array_1509 AND_array_1509_c615({a_c[893:0],615'd0},p_prime[615],c_w_615);
AND_array_1509 AND_array_1509_s615({a_s[893:0],615'd0},p_prime[615],s_w_615);
AND_array_1509 AND_array_1509_c616({a_c[892:0],616'd0},p_prime[616],c_w_616);
AND_array_1509 AND_array_1509_s616({a_s[892:0],616'd0},p_prime[616],s_w_616);
AND_array_1509 AND_array_1509_c617({a_c[891:0],617'd0},p_prime[617],c_w_617);
AND_array_1509 AND_array_1509_s617({a_s[891:0],617'd0},p_prime[617],s_w_617);
AND_array_1509 AND_array_1509_c618({a_c[890:0],618'd0},p_prime[618],c_w_618);
AND_array_1509 AND_array_1509_s618({a_s[890:0],618'd0},p_prime[618],s_w_618);
AND_array_1509 AND_array_1509_c619({a_c[889:0],619'd0},p_prime[619],c_w_619);
AND_array_1509 AND_array_1509_s619({a_s[889:0],619'd0},p_prime[619],s_w_619);
AND_array_1509 AND_array_1509_c620({a_c[888:0],620'd0},p_prime[620],c_w_620);
AND_array_1509 AND_array_1509_s620({a_s[888:0],620'd0},p_prime[620],s_w_620);
AND_array_1509 AND_array_1509_c621({a_c[887:0],621'd0},p_prime[621],c_w_621);
AND_array_1509 AND_array_1509_s621({a_s[887:0],621'd0},p_prime[621],s_w_621);
AND_array_1509 AND_array_1509_c622({a_c[886:0],622'd0},p_prime[622],c_w_622);
AND_array_1509 AND_array_1509_s622({a_s[886:0],622'd0},p_prime[622],s_w_622);
AND_array_1509 AND_array_1509_c623({a_c[885:0],623'd0},p_prime[623],c_w_623);
AND_array_1509 AND_array_1509_s623({a_s[885:0],623'd0},p_prime[623],s_w_623);
AND_array_1509 AND_array_1509_c624({a_c[884:0],624'd0},p_prime[624],c_w_624);
AND_array_1509 AND_array_1509_s624({a_s[884:0],624'd0},p_prime[624],s_w_624);
AND_array_1509 AND_array_1509_c625({a_c[883:0],625'd0},p_prime[625],c_w_625);
AND_array_1509 AND_array_1509_s625({a_s[883:0],625'd0},p_prime[625],s_w_625);
AND_array_1509 AND_array_1509_c626({a_c[882:0],626'd0},p_prime[626],c_w_626);
AND_array_1509 AND_array_1509_s626({a_s[882:0],626'd0},p_prime[626],s_w_626);
AND_array_1509 AND_array_1509_c627({a_c[881:0],627'd0},p_prime[627],c_w_627);
AND_array_1509 AND_array_1509_s627({a_s[881:0],627'd0},p_prime[627],s_w_627);
AND_array_1509 AND_array_1509_c628({a_c[880:0],628'd0},p_prime[628],c_w_628);
AND_array_1509 AND_array_1509_s628({a_s[880:0],628'd0},p_prime[628],s_w_628);
AND_array_1509 AND_array_1509_c629({a_c[879:0],629'd0},p_prime[629],c_w_629);
AND_array_1509 AND_array_1509_s629({a_s[879:0],629'd0},p_prime[629],s_w_629);
AND_array_1509 AND_array_1509_c630({a_c[878:0],630'd0},p_prime[630],c_w_630);
AND_array_1509 AND_array_1509_s630({a_s[878:0],630'd0},p_prime[630],s_w_630);
AND_array_1509 AND_array_1509_c631({a_c[877:0],631'd0},p_prime[631],c_w_631);
AND_array_1509 AND_array_1509_s631({a_s[877:0],631'd0},p_prime[631],s_w_631);
AND_array_1509 AND_array_1509_c632({a_c[876:0],632'd0},p_prime[632],c_w_632);
AND_array_1509 AND_array_1509_s632({a_s[876:0],632'd0},p_prime[632],s_w_632);
AND_array_1509 AND_array_1509_c633({a_c[875:0],633'd0},p_prime[633],c_w_633);
AND_array_1509 AND_array_1509_s633({a_s[875:0],633'd0},p_prime[633],s_w_633);
AND_array_1509 AND_array_1509_c634({a_c[874:0],634'd0},p_prime[634],c_w_634);
AND_array_1509 AND_array_1509_s634({a_s[874:0],634'd0},p_prime[634],s_w_634);
AND_array_1509 AND_array_1509_c635({a_c[873:0],635'd0},p_prime[635],c_w_635);
AND_array_1509 AND_array_1509_s635({a_s[873:0],635'd0},p_prime[635],s_w_635);
AND_array_1509 AND_array_1509_c636({a_c[872:0],636'd0},p_prime[636],c_w_636);
AND_array_1509 AND_array_1509_s636({a_s[872:0],636'd0},p_prime[636],s_w_636);
AND_array_1509 AND_array_1509_c637({a_c[871:0],637'd0},p_prime[637],c_w_637);
AND_array_1509 AND_array_1509_s637({a_s[871:0],637'd0},p_prime[637],s_w_637);
AND_array_1509 AND_array_1509_c638({a_c[870:0],638'd0},p_prime[638],c_w_638);
AND_array_1509 AND_array_1509_s638({a_s[870:0],638'd0},p_prime[638],s_w_638);
AND_array_1509 AND_array_1509_c639({a_c[869:0],639'd0},p_prime[639],c_w_639);
AND_array_1509 AND_array_1509_s639({a_s[869:0],639'd0},p_prime[639],s_w_639);
AND_array_1509 AND_array_1509_c640({a_c[868:0],640'd0},p_prime[640],c_w_640);
AND_array_1509 AND_array_1509_s640({a_s[868:0],640'd0},p_prime[640],s_w_640);
AND_array_1509 AND_array_1509_c641({a_c[867:0],641'd0},p_prime[641],c_w_641);
AND_array_1509 AND_array_1509_s641({a_s[867:0],641'd0},p_prime[641],s_w_641);
AND_array_1509 AND_array_1509_c642({a_c[866:0],642'd0},p_prime[642],c_w_642);
AND_array_1509 AND_array_1509_s642({a_s[866:0],642'd0},p_prime[642],s_w_642);
AND_array_1509 AND_array_1509_c643({a_c[865:0],643'd0},p_prime[643],c_w_643);
AND_array_1509 AND_array_1509_s643({a_s[865:0],643'd0},p_prime[643],s_w_643);
AND_array_1509 AND_array_1509_c644({a_c[864:0],644'd0},p_prime[644],c_w_644);
AND_array_1509 AND_array_1509_s644({a_s[864:0],644'd0},p_prime[644],s_w_644);
AND_array_1509 AND_array_1509_c645({a_c[863:0],645'd0},p_prime[645],c_w_645);
AND_array_1509 AND_array_1509_s645({a_s[863:0],645'd0},p_prime[645],s_w_645);
AND_array_1509 AND_array_1509_c646({a_c[862:0],646'd0},p_prime[646],c_w_646);
AND_array_1509 AND_array_1509_s646({a_s[862:0],646'd0},p_prime[646],s_w_646);
AND_array_1509 AND_array_1509_c647({a_c[861:0],647'd0},p_prime[647],c_w_647);
AND_array_1509 AND_array_1509_s647({a_s[861:0],647'd0},p_prime[647],s_w_647);
AND_array_1509 AND_array_1509_c648({a_c[860:0],648'd0},p_prime[648],c_w_648);
AND_array_1509 AND_array_1509_s648({a_s[860:0],648'd0},p_prime[648],s_w_648);
AND_array_1509 AND_array_1509_c649({a_c[859:0],649'd0},p_prime[649],c_w_649);
AND_array_1509 AND_array_1509_s649({a_s[859:0],649'd0},p_prime[649],s_w_649);
AND_array_1509 AND_array_1509_c650({a_c[858:0],650'd0},p_prime[650],c_w_650);
AND_array_1509 AND_array_1509_s650({a_s[858:0],650'd0},p_prime[650],s_w_650);
AND_array_1509 AND_array_1509_c651({a_c[857:0],651'd0},p_prime[651],c_w_651);
AND_array_1509 AND_array_1509_s651({a_s[857:0],651'd0},p_prime[651],s_w_651);
AND_array_1509 AND_array_1509_c652({a_c[856:0],652'd0},p_prime[652],c_w_652);
AND_array_1509 AND_array_1509_s652({a_s[856:0],652'd0},p_prime[652],s_w_652);
AND_array_1509 AND_array_1509_c653({a_c[855:0],653'd0},p_prime[653],c_w_653);
AND_array_1509 AND_array_1509_s653({a_s[855:0],653'd0},p_prime[653],s_w_653);
AND_array_1509 AND_array_1509_c654({a_c[854:0],654'd0},p_prime[654],c_w_654);
AND_array_1509 AND_array_1509_s654({a_s[854:0],654'd0},p_prime[654],s_w_654);
AND_array_1509 AND_array_1509_c655({a_c[853:0],655'd0},p_prime[655],c_w_655);
AND_array_1509 AND_array_1509_s655({a_s[853:0],655'd0},p_prime[655],s_w_655);
AND_array_1509 AND_array_1509_c656({a_c[852:0],656'd0},p_prime[656],c_w_656);
AND_array_1509 AND_array_1509_s656({a_s[852:0],656'd0},p_prime[656],s_w_656);
AND_array_1509 AND_array_1509_c657({a_c[851:0],657'd0},p_prime[657],c_w_657);
AND_array_1509 AND_array_1509_s657({a_s[851:0],657'd0},p_prime[657],s_w_657);
AND_array_1509 AND_array_1509_c658({a_c[850:0],658'd0},p_prime[658],c_w_658);
AND_array_1509 AND_array_1509_s658({a_s[850:0],658'd0},p_prime[658],s_w_658);
AND_array_1509 AND_array_1509_c659({a_c[849:0],659'd0},p_prime[659],c_w_659);
AND_array_1509 AND_array_1509_s659({a_s[849:0],659'd0},p_prime[659],s_w_659);
AND_array_1509 AND_array_1509_c660({a_c[848:0],660'd0},p_prime[660],c_w_660);
AND_array_1509 AND_array_1509_s660({a_s[848:0],660'd0},p_prime[660],s_w_660);
AND_array_1509 AND_array_1509_c661({a_c[847:0],661'd0},p_prime[661],c_w_661);
AND_array_1509 AND_array_1509_s661({a_s[847:0],661'd0},p_prime[661],s_w_661);
AND_array_1509 AND_array_1509_c662({a_c[846:0],662'd0},p_prime[662],c_w_662);
AND_array_1509 AND_array_1509_s662({a_s[846:0],662'd0},p_prime[662],s_w_662);
AND_array_1509 AND_array_1509_c663({a_c[845:0],663'd0},p_prime[663],c_w_663);
AND_array_1509 AND_array_1509_s663({a_s[845:0],663'd0},p_prime[663],s_w_663);
AND_array_1509 AND_array_1509_c664({a_c[844:0],664'd0},p_prime[664],c_w_664);
AND_array_1509 AND_array_1509_s664({a_s[844:0],664'd0},p_prime[664],s_w_664);
AND_array_1509 AND_array_1509_c665({a_c[843:0],665'd0},p_prime[665],c_w_665);
AND_array_1509 AND_array_1509_s665({a_s[843:0],665'd0},p_prime[665],s_w_665);
AND_array_1509 AND_array_1509_c666({a_c[842:0],666'd0},p_prime[666],c_w_666);
AND_array_1509 AND_array_1509_s666({a_s[842:0],666'd0},p_prime[666],s_w_666);
AND_array_1509 AND_array_1509_c667({a_c[841:0],667'd0},p_prime[667],c_w_667);
AND_array_1509 AND_array_1509_s667({a_s[841:0],667'd0},p_prime[667],s_w_667);
AND_array_1509 AND_array_1509_c668({a_c[840:0],668'd0},p_prime[668],c_w_668);
AND_array_1509 AND_array_1509_s668({a_s[840:0],668'd0},p_prime[668],s_w_668);
AND_array_1509 AND_array_1509_c669({a_c[839:0],669'd0},p_prime[669],c_w_669);
AND_array_1509 AND_array_1509_s669({a_s[839:0],669'd0},p_prime[669],s_w_669);
AND_array_1509 AND_array_1509_c670({a_c[838:0],670'd0},p_prime[670],c_w_670);
AND_array_1509 AND_array_1509_s670({a_s[838:0],670'd0},p_prime[670],s_w_670);
AND_array_1509 AND_array_1509_c671({a_c[837:0],671'd0},p_prime[671],c_w_671);
AND_array_1509 AND_array_1509_s671({a_s[837:0],671'd0},p_prime[671],s_w_671);
AND_array_1509 AND_array_1509_c672({a_c[836:0],672'd0},p_prime[672],c_w_672);
AND_array_1509 AND_array_1509_s672({a_s[836:0],672'd0},p_prime[672],s_w_672);
AND_array_1509 AND_array_1509_c673({a_c[835:0],673'd0},p_prime[673],c_w_673);
AND_array_1509 AND_array_1509_s673({a_s[835:0],673'd0},p_prime[673],s_w_673);
AND_array_1509 AND_array_1509_c674({a_c[834:0],674'd0},p_prime[674],c_w_674);
AND_array_1509 AND_array_1509_s674({a_s[834:0],674'd0},p_prime[674],s_w_674);
AND_array_1509 AND_array_1509_c675({a_c[833:0],675'd0},p_prime[675],c_w_675);
AND_array_1509 AND_array_1509_s675({a_s[833:0],675'd0},p_prime[675],s_w_675);
AND_array_1509 AND_array_1509_c676({a_c[832:0],676'd0},p_prime[676],c_w_676);
AND_array_1509 AND_array_1509_s676({a_s[832:0],676'd0},p_prime[676],s_w_676);
AND_array_1509 AND_array_1509_c677({a_c[831:0],677'd0},p_prime[677],c_w_677);
AND_array_1509 AND_array_1509_s677({a_s[831:0],677'd0},p_prime[677],s_w_677);
AND_array_1509 AND_array_1509_c678({a_c[830:0],678'd0},p_prime[678],c_w_678);
AND_array_1509 AND_array_1509_s678({a_s[830:0],678'd0},p_prime[678],s_w_678);
AND_array_1509 AND_array_1509_c679({a_c[829:0],679'd0},p_prime[679],c_w_679);
AND_array_1509 AND_array_1509_s679({a_s[829:0],679'd0},p_prime[679],s_w_679);
AND_array_1509 AND_array_1509_c680({a_c[828:0],680'd0},p_prime[680],c_w_680);
AND_array_1509 AND_array_1509_s680({a_s[828:0],680'd0},p_prime[680],s_w_680);
AND_array_1509 AND_array_1509_c681({a_c[827:0],681'd0},p_prime[681],c_w_681);
AND_array_1509 AND_array_1509_s681({a_s[827:0],681'd0},p_prime[681],s_w_681);
AND_array_1509 AND_array_1509_c682({a_c[826:0],682'd0},p_prime[682],c_w_682);
AND_array_1509 AND_array_1509_s682({a_s[826:0],682'd0},p_prime[682],s_w_682);
AND_array_1509 AND_array_1509_c683({a_c[825:0],683'd0},p_prime[683],c_w_683);
AND_array_1509 AND_array_1509_s683({a_s[825:0],683'd0},p_prime[683],s_w_683);
AND_array_1509 AND_array_1509_c684({a_c[824:0],684'd0},p_prime[684],c_w_684);
AND_array_1509 AND_array_1509_s684({a_s[824:0],684'd0},p_prime[684],s_w_684);
AND_array_1509 AND_array_1509_c685({a_c[823:0],685'd0},p_prime[685],c_w_685);
AND_array_1509 AND_array_1509_s685({a_s[823:0],685'd0},p_prime[685],s_w_685);
AND_array_1509 AND_array_1509_c686({a_c[822:0],686'd0},p_prime[686],c_w_686);
AND_array_1509 AND_array_1509_s686({a_s[822:0],686'd0},p_prime[686],s_w_686);
AND_array_1509 AND_array_1509_c687({a_c[821:0],687'd0},p_prime[687],c_w_687);
AND_array_1509 AND_array_1509_s687({a_s[821:0],687'd0},p_prime[687],s_w_687);
AND_array_1509 AND_array_1509_c688({a_c[820:0],688'd0},p_prime[688],c_w_688);
AND_array_1509 AND_array_1509_s688({a_s[820:0],688'd0},p_prime[688],s_w_688);
AND_array_1509 AND_array_1509_c689({a_c[819:0],689'd0},p_prime[689],c_w_689);
AND_array_1509 AND_array_1509_s689({a_s[819:0],689'd0},p_prime[689],s_w_689);
AND_array_1509 AND_array_1509_c690({a_c[818:0],690'd0},p_prime[690],c_w_690);
AND_array_1509 AND_array_1509_s690({a_s[818:0],690'd0},p_prime[690],s_w_690);
AND_array_1509 AND_array_1509_c691({a_c[817:0],691'd0},p_prime[691],c_w_691);
AND_array_1509 AND_array_1509_s691({a_s[817:0],691'd0},p_prime[691],s_w_691);
AND_array_1509 AND_array_1509_c692({a_c[816:0],692'd0},p_prime[692],c_w_692);
AND_array_1509 AND_array_1509_s692({a_s[816:0],692'd0},p_prime[692],s_w_692);
AND_array_1509 AND_array_1509_c693({a_c[815:0],693'd0},p_prime[693],c_w_693);
AND_array_1509 AND_array_1509_s693({a_s[815:0],693'd0},p_prime[693],s_w_693);
AND_array_1509 AND_array_1509_c694({a_c[814:0],694'd0},p_prime[694],c_w_694);
AND_array_1509 AND_array_1509_s694({a_s[814:0],694'd0},p_prime[694],s_w_694);
AND_array_1509 AND_array_1509_c695({a_c[813:0],695'd0},p_prime[695],c_w_695);
AND_array_1509 AND_array_1509_s695({a_s[813:0],695'd0},p_prime[695],s_w_695);
AND_array_1509 AND_array_1509_c696({a_c[812:0],696'd0},p_prime[696],c_w_696);
AND_array_1509 AND_array_1509_s696({a_s[812:0],696'd0},p_prime[696],s_w_696);
AND_array_1509 AND_array_1509_c697({a_c[811:0],697'd0},p_prime[697],c_w_697);
AND_array_1509 AND_array_1509_s697({a_s[811:0],697'd0},p_prime[697],s_w_697);
AND_array_1509 AND_array_1509_c698({a_c[810:0],698'd0},p_prime[698],c_w_698);
AND_array_1509 AND_array_1509_s698({a_s[810:0],698'd0},p_prime[698],s_w_698);
AND_array_1509 AND_array_1509_c699({a_c[809:0],699'd0},p_prime[699],c_w_699);
AND_array_1509 AND_array_1509_s699({a_s[809:0],699'd0},p_prime[699],s_w_699);
AND_array_1509 AND_array_1509_c700({a_c[808:0],700'd0},p_prime[700],c_w_700);
AND_array_1509 AND_array_1509_s700({a_s[808:0],700'd0},p_prime[700],s_w_700);
AND_array_1509 AND_array_1509_c701({a_c[807:0],701'd0},p_prime[701],c_w_701);
AND_array_1509 AND_array_1509_s701({a_s[807:0],701'd0},p_prime[701],s_w_701);
AND_array_1509 AND_array_1509_c702({a_c[806:0],702'd0},p_prime[702],c_w_702);
AND_array_1509 AND_array_1509_s702({a_s[806:0],702'd0},p_prime[702],s_w_702);
AND_array_1509 AND_array_1509_c703({a_c[805:0],703'd0},p_prime[703],c_w_703);
AND_array_1509 AND_array_1509_s703({a_s[805:0],703'd0},p_prime[703],s_w_703);
AND_array_1509 AND_array_1509_c704({a_c[804:0],704'd0},p_prime[704],c_w_704);
AND_array_1509 AND_array_1509_s704({a_s[804:0],704'd0},p_prime[704],s_w_704);
AND_array_1509 AND_array_1509_c705({a_c[803:0],705'd0},p_prime[705],c_w_705);
AND_array_1509 AND_array_1509_s705({a_s[803:0],705'd0},p_prime[705],s_w_705);
AND_array_1509 AND_array_1509_c706({a_c[802:0],706'd0},p_prime[706],c_w_706);
AND_array_1509 AND_array_1509_s706({a_s[802:0],706'd0},p_prime[706],s_w_706);
AND_array_1509 AND_array_1509_c707({a_c[801:0],707'd0},p_prime[707],c_w_707);
AND_array_1509 AND_array_1509_s707({a_s[801:0],707'd0},p_prime[707],s_w_707);
AND_array_1509 AND_array_1509_c708({a_c[800:0],708'd0},p_prime[708],c_w_708);
AND_array_1509 AND_array_1509_s708({a_s[800:0],708'd0},p_prime[708],s_w_708);
AND_array_1509 AND_array_1509_c709({a_c[799:0],709'd0},p_prime[709],c_w_709);
AND_array_1509 AND_array_1509_s709({a_s[799:0],709'd0},p_prime[709],s_w_709);
AND_array_1509 AND_array_1509_c710({a_c[798:0],710'd0},p_prime[710],c_w_710);
AND_array_1509 AND_array_1509_s710({a_s[798:0],710'd0},p_prime[710],s_w_710);
AND_array_1509 AND_array_1509_c711({a_c[797:0],711'd0},p_prime[711],c_w_711);
AND_array_1509 AND_array_1509_s711({a_s[797:0],711'd0},p_prime[711],s_w_711);
AND_array_1509 AND_array_1509_c712({a_c[796:0],712'd0},p_prime[712],c_w_712);
AND_array_1509 AND_array_1509_s712({a_s[796:0],712'd0},p_prime[712],s_w_712);
AND_array_1509 AND_array_1509_c713({a_c[795:0],713'd0},p_prime[713],c_w_713);
AND_array_1509 AND_array_1509_s713({a_s[795:0],713'd0},p_prime[713],s_w_713);
AND_array_1509 AND_array_1509_c714({a_c[794:0],714'd0},p_prime[714],c_w_714);
AND_array_1509 AND_array_1509_s714({a_s[794:0],714'd0},p_prime[714],s_w_714);
AND_array_1509 AND_array_1509_c715({a_c[793:0],715'd0},p_prime[715],c_w_715);
AND_array_1509 AND_array_1509_s715({a_s[793:0],715'd0},p_prime[715],s_w_715);
AND_array_1509 AND_array_1509_c716({a_c[792:0],716'd0},p_prime[716],c_w_716);
AND_array_1509 AND_array_1509_s716({a_s[792:0],716'd0},p_prime[716],s_w_716);
AND_array_1509 AND_array_1509_c717({a_c[791:0],717'd0},p_prime[717],c_w_717);
AND_array_1509 AND_array_1509_s717({a_s[791:0],717'd0},p_prime[717],s_w_717);
AND_array_1509 AND_array_1509_c718({a_c[790:0],718'd0},p_prime[718],c_w_718);
AND_array_1509 AND_array_1509_s718({a_s[790:0],718'd0},p_prime[718],s_w_718);
AND_array_1509 AND_array_1509_c719({a_c[789:0],719'd0},p_prime[719],c_w_719);
AND_array_1509 AND_array_1509_s719({a_s[789:0],719'd0},p_prime[719],s_w_719);
AND_array_1509 AND_array_1509_c720({a_c[788:0],720'd0},p_prime[720],c_w_720);
AND_array_1509 AND_array_1509_s720({a_s[788:0],720'd0},p_prime[720],s_w_720);
AND_array_1509 AND_array_1509_c721({a_c[787:0],721'd0},p_prime[721],c_w_721);
AND_array_1509 AND_array_1509_s721({a_s[787:0],721'd0},p_prime[721],s_w_721);
AND_array_1509 AND_array_1509_c722({a_c[786:0],722'd0},p_prime[722],c_w_722);
AND_array_1509 AND_array_1509_s722({a_s[786:0],722'd0},p_prime[722],s_w_722);
AND_array_1509 AND_array_1509_c723({a_c[785:0],723'd0},p_prime[723],c_w_723);
AND_array_1509 AND_array_1509_s723({a_s[785:0],723'd0},p_prime[723],s_w_723);
AND_array_1509 AND_array_1509_c724({a_c[784:0],724'd0},p_prime[724],c_w_724);
AND_array_1509 AND_array_1509_s724({a_s[784:0],724'd0},p_prime[724],s_w_724);
AND_array_1509 AND_array_1509_c725({a_c[783:0],725'd0},p_prime[725],c_w_725);
AND_array_1509 AND_array_1509_s725({a_s[783:0],725'd0},p_prime[725],s_w_725);
AND_array_1509 AND_array_1509_c726({a_c[782:0],726'd0},p_prime[726],c_w_726);
AND_array_1509 AND_array_1509_s726({a_s[782:0],726'd0},p_prime[726],s_w_726);
AND_array_1509 AND_array_1509_c727({a_c[781:0],727'd0},p_prime[727],c_w_727);
AND_array_1509 AND_array_1509_s727({a_s[781:0],727'd0},p_prime[727],s_w_727);
AND_array_1509 AND_array_1509_c728({a_c[780:0],728'd0},p_prime[728],c_w_728);
AND_array_1509 AND_array_1509_s728({a_s[780:0],728'd0},p_prime[728],s_w_728);
AND_array_1509 AND_array_1509_c729({a_c[779:0],729'd0},p_prime[729],c_w_729);
AND_array_1509 AND_array_1509_s729({a_s[779:0],729'd0},p_prime[729],s_w_729);
AND_array_1509 AND_array_1509_c730({a_c[778:0],730'd0},p_prime[730],c_w_730);
AND_array_1509 AND_array_1509_s730({a_s[778:0],730'd0},p_prime[730],s_w_730);
AND_array_1509 AND_array_1509_c731({a_c[777:0],731'd0},p_prime[731],c_w_731);
AND_array_1509 AND_array_1509_s731({a_s[777:0],731'd0},p_prime[731],s_w_731);
AND_array_1509 AND_array_1509_c732({a_c[776:0],732'd0},p_prime[732],c_w_732);
AND_array_1509 AND_array_1509_s732({a_s[776:0],732'd0},p_prime[732],s_w_732);
AND_array_1509 AND_array_1509_c733({a_c[775:0],733'd0},p_prime[733],c_w_733);
AND_array_1509 AND_array_1509_s733({a_s[775:0],733'd0},p_prime[733],s_w_733);
AND_array_1509 AND_array_1509_c734({a_c[774:0],734'd0},p_prime[734],c_w_734);
AND_array_1509 AND_array_1509_s734({a_s[774:0],734'd0},p_prime[734],s_w_734);
AND_array_1509 AND_array_1509_c735({a_c[773:0],735'd0},p_prime[735],c_w_735);
AND_array_1509 AND_array_1509_s735({a_s[773:0],735'd0},p_prime[735],s_w_735);
AND_array_1509 AND_array_1509_c736({a_c[772:0],736'd0},p_prime[736],c_w_736);
AND_array_1509 AND_array_1509_s736({a_s[772:0],736'd0},p_prime[736],s_w_736);
AND_array_1509 AND_array_1509_c737({a_c[771:0],737'd0},p_prime[737],c_w_737);
AND_array_1509 AND_array_1509_s737({a_s[771:0],737'd0},p_prime[737],s_w_737);
AND_array_1509 AND_array_1509_c738({a_c[770:0],738'd0},p_prime[738],c_w_738);
AND_array_1509 AND_array_1509_s738({a_s[770:0],738'd0},p_prime[738],s_w_738);
AND_array_1509 AND_array_1509_c739({a_c[769:0],739'd0},p_prime[739],c_w_739);
AND_array_1509 AND_array_1509_s739({a_s[769:0],739'd0},p_prime[739],s_w_739);
AND_array_1509 AND_array_1509_c740({a_c[768:0],740'd0},p_prime[740],c_w_740);
AND_array_1509 AND_array_1509_s740({a_s[768:0],740'd0},p_prime[740],s_w_740);
AND_array_1509 AND_array_1509_c741({a_c[767:0],741'd0},p_prime[741],c_w_741);
AND_array_1509 AND_array_1509_s741({a_s[767:0],741'd0},p_prime[741],s_w_741);
AND_array_1509 AND_array_1509_c742({a_c[766:0],742'd0},p_prime[742],c_w_742);
AND_array_1509 AND_array_1509_s742({a_s[766:0],742'd0},p_prime[742],s_w_742);
AND_array_1509 AND_array_1509_c743({a_c[765:0],743'd0},p_prime[743],c_w_743);
AND_array_1509 AND_array_1509_s743({a_s[765:0],743'd0},p_prime[743],s_w_743);
AND_array_1509 AND_array_1509_c744({a_c[764:0],744'd0},p_prime[744],c_w_744);
AND_array_1509 AND_array_1509_s744({a_s[764:0],744'd0},p_prime[744],s_w_744);
AND_array_1509 AND_array_1509_c745({a_c[763:0],745'd0},p_prime[745],c_w_745);
AND_array_1509 AND_array_1509_s745({a_s[763:0],745'd0},p_prime[745],s_w_745);
AND_array_1509 AND_array_1509_c746({a_c[762:0],746'd0},p_prime[746],c_w_746);
AND_array_1509 AND_array_1509_s746({a_s[762:0],746'd0},p_prime[746],s_w_746);
AND_array_1509 AND_array_1509_c747({a_c[761:0],747'd0},p_prime[747],c_w_747);
AND_array_1509 AND_array_1509_s747({a_s[761:0],747'd0},p_prime[747],s_w_747);
AND_array_1509 AND_array_1509_c748({a_c[760:0],748'd0},p_prime[748],c_w_748);
AND_array_1509 AND_array_1509_s748({a_s[760:0],748'd0},p_prime[748],s_w_748);
AND_array_1509 AND_array_1509_c749({a_c[759:0],749'd0},p_prime[749],c_w_749);
AND_array_1509 AND_array_1509_s749({a_s[759:0],749'd0},p_prime[749],s_w_749);
AND_array_1509 AND_array_1509_c750({a_c[758:0],750'd0},p_prime[750],c_w_750);
AND_array_1509 AND_array_1509_s750({a_s[758:0],750'd0},p_prime[750],s_w_750);
AND_array_1509 AND_array_1509_c751({a_c[757:0],751'd0},p_prime[751],c_w_751);
AND_array_1509 AND_array_1509_s751({a_s[757:0],751'd0},p_prime[751],s_w_751);
AND_array_1509 AND_array_1509_c752({a_c[756:0],752'd0},p_prime[752],c_w_752);
AND_array_1509 AND_array_1509_s752({a_s[756:0],752'd0},p_prime[752],s_w_752);
AND_array_1509 AND_array_1509_c753({a_c[755:0],753'd0},p_prime[753],c_w_753);
AND_array_1509 AND_array_1509_s753({a_s[755:0],753'd0},p_prime[753],s_w_753);
AND_array_1509 AND_array_1509_c754({a_c[754:0],754'd0},p_prime[754],c_w_754);
AND_array_1509 AND_array_1509_s754({a_s[754:0],754'd0},p_prime[754],s_w_754);
AND_array_1509 AND_array_1509_c755({a_c[753:0],755'd0},p_prime[755],c_w_755);
AND_array_1509 AND_array_1509_s755({a_s[753:0],755'd0},p_prime[755],s_w_755);
AND_array_1509 AND_array_1509_c756({a_c[752:0],756'd0},p_prime[756],c_w_756);
AND_array_1509 AND_array_1509_s756({a_s[752:0],756'd0},p_prime[756],s_w_756);
AND_array_1509 AND_array_1509_c757({a_c[751:0],757'd0},p_prime[757],c_w_757);
AND_array_1509 AND_array_1509_s757({a_s[751:0],757'd0},p_prime[757],s_w_757);
AND_array_1509 AND_array_1509_c758({a_c[750:0],758'd0},p_prime[758],c_w_758);
AND_array_1509 AND_array_1509_s758({a_s[750:0],758'd0},p_prime[758],s_w_758);
AND_array_1509 AND_array_1509_c759({a_c[749:0],759'd0},p_prime[759],c_w_759);
AND_array_1509 AND_array_1509_s759({a_s[749:0],759'd0},p_prime[759],s_w_759);
AND_array_1509 AND_array_1509_c760({a_c[748:0],760'd0},p_prime[760],c_w_760);
AND_array_1509 AND_array_1509_s760({a_s[748:0],760'd0},p_prime[760],s_w_760);
AND_array_1509 AND_array_1509_c761({a_c[747:0],761'd0},p_prime[761],c_w_761);
AND_array_1509 AND_array_1509_s761({a_s[747:0],761'd0},p_prime[761],s_w_761);
AND_array_1509 AND_array_1509_c762({a_c[746:0],762'd0},p_prime[762],c_w_762);
AND_array_1509 AND_array_1509_s762({a_s[746:0],762'd0},p_prime[762],s_w_762);
AND_array_1509 AND_array_1509_c763({a_c[745:0],763'd0},p_prime[763],c_w_763);
AND_array_1509 AND_array_1509_s763({a_s[745:0],763'd0},p_prime[763],s_w_763);
AND_array_1509 AND_array_1509_c764({a_c[744:0],764'd0},p_prime[764],c_w_764);
AND_array_1509 AND_array_1509_s764({a_s[744:0],764'd0},p_prime[764],s_w_764);
AND_array_1509 AND_array_1509_c765({a_c[743:0],765'd0},p_prime[765],c_w_765);
AND_array_1509 AND_array_1509_s765({a_s[743:0],765'd0},p_prime[765],s_w_765);
AND_array_1509 AND_array_1509_c766({a_c[742:0],766'd0},p_prime[766],c_w_766);
AND_array_1509 AND_array_1509_s766({a_s[742:0],766'd0},p_prime[766],s_w_766);
AND_array_1509 AND_array_1509_c767({a_c[741:0],767'd0},p_prime[767],c_w_767);
AND_array_1509 AND_array_1509_s767({a_s[741:0],767'd0},p_prime[767],s_w_767);
AND_array_1509 AND_array_1509_c768({a_c[740:0],768'd0},p_prime[768],c_w_768);
AND_array_1509 AND_array_1509_s768({a_s[740:0],768'd0},p_prime[768],s_w_768);
AND_array_1509 AND_array_1509_c769({a_c[739:0],769'd0},p_prime[769],c_w_769);
AND_array_1509 AND_array_1509_s769({a_s[739:0],769'd0},p_prime[769],s_w_769);
AND_array_1509 AND_array_1509_c770({a_c[738:0],770'd0},p_prime[770],c_w_770);
AND_array_1509 AND_array_1509_s770({a_s[738:0],770'd0},p_prime[770],s_w_770);
AND_array_1509 AND_array_1509_c771({a_c[737:0],771'd0},p_prime[771],c_w_771);
AND_array_1509 AND_array_1509_s771({a_s[737:0],771'd0},p_prime[771],s_w_771);
AND_array_1509 AND_array_1509_c772({a_c[736:0],772'd0},p_prime[772],c_w_772);
AND_array_1509 AND_array_1509_s772({a_s[736:0],772'd0},p_prime[772],s_w_772);
AND_array_1509 AND_array_1509_c773({a_c[735:0],773'd0},p_prime[773],c_w_773);
AND_array_1509 AND_array_1509_s773({a_s[735:0],773'd0},p_prime[773],s_w_773);
AND_array_1509 AND_array_1509_c774({a_c[734:0],774'd0},p_prime[774],c_w_774);
AND_array_1509 AND_array_1509_s774({a_s[734:0],774'd0},p_prime[774],s_w_774);
AND_array_1509 AND_array_1509_c775({a_c[733:0],775'd0},p_prime[775],c_w_775);
AND_array_1509 AND_array_1509_s775({a_s[733:0],775'd0},p_prime[775],s_w_775);
AND_array_1509 AND_array_1509_c776({a_c[732:0],776'd0},p_prime[776],c_w_776);
AND_array_1509 AND_array_1509_s776({a_s[732:0],776'd0},p_prime[776],s_w_776);
AND_array_1509 AND_array_1509_c777({a_c[731:0],777'd0},p_prime[777],c_w_777);
AND_array_1509 AND_array_1509_s777({a_s[731:0],777'd0},p_prime[777],s_w_777);
AND_array_1509 AND_array_1509_c778({a_c[730:0],778'd0},p_prime[778],c_w_778);
AND_array_1509 AND_array_1509_s778({a_s[730:0],778'd0},p_prime[778],s_w_778);
AND_array_1509 AND_array_1509_c779({a_c[729:0],779'd0},p_prime[779],c_w_779);
AND_array_1509 AND_array_1509_s779({a_s[729:0],779'd0},p_prime[779],s_w_779);
AND_array_1509 AND_array_1509_c780({a_c[728:0],780'd0},p_prime[780],c_w_780);
AND_array_1509 AND_array_1509_s780({a_s[728:0],780'd0},p_prime[780],s_w_780);
AND_array_1509 AND_array_1509_c781({a_c[727:0],781'd0},p_prime[781],c_w_781);
AND_array_1509 AND_array_1509_s781({a_s[727:0],781'd0},p_prime[781],s_w_781);
AND_array_1509 AND_array_1509_c782({a_c[726:0],782'd0},p_prime[782],c_w_782);
AND_array_1509 AND_array_1509_s782({a_s[726:0],782'd0},p_prime[782],s_w_782);
AND_array_1509 AND_array_1509_c783({a_c[725:0],783'd0},p_prime[783],c_w_783);
AND_array_1509 AND_array_1509_s783({a_s[725:0],783'd0},p_prime[783],s_w_783);
AND_array_1509 AND_array_1509_c784({a_c[724:0],784'd0},p_prime[784],c_w_784);
AND_array_1509 AND_array_1509_s784({a_s[724:0],784'd0},p_prime[784],s_w_784);
AND_array_1509 AND_array_1509_c785({a_c[723:0],785'd0},p_prime[785],c_w_785);
AND_array_1509 AND_array_1509_s785({a_s[723:0],785'd0},p_prime[785],s_w_785);
AND_array_1509 AND_array_1509_c786({a_c[722:0],786'd0},p_prime[786],c_w_786);
AND_array_1509 AND_array_1509_s786({a_s[722:0],786'd0},p_prime[786],s_w_786);
AND_array_1509 AND_array_1509_c787({a_c[721:0],787'd0},p_prime[787],c_w_787);
AND_array_1509 AND_array_1509_s787({a_s[721:0],787'd0},p_prime[787],s_w_787);
AND_array_1509 AND_array_1509_c788({a_c[720:0],788'd0},p_prime[788],c_w_788);
AND_array_1509 AND_array_1509_s788({a_s[720:0],788'd0},p_prime[788],s_w_788);
AND_array_1509 AND_array_1509_c789({a_c[719:0],789'd0},p_prime[789],c_w_789);
AND_array_1509 AND_array_1509_s789({a_s[719:0],789'd0},p_prime[789],s_w_789);
AND_array_1509 AND_array_1509_c790({a_c[718:0],790'd0},p_prime[790],c_w_790);
AND_array_1509 AND_array_1509_s790({a_s[718:0],790'd0},p_prime[790],s_w_790);
AND_array_1509 AND_array_1509_c791({a_c[717:0],791'd0},p_prime[791],c_w_791);
AND_array_1509 AND_array_1509_s791({a_s[717:0],791'd0},p_prime[791],s_w_791);
AND_array_1509 AND_array_1509_c792({a_c[716:0],792'd0},p_prime[792],c_w_792);
AND_array_1509 AND_array_1509_s792({a_s[716:0],792'd0},p_prime[792],s_w_792);
AND_array_1509 AND_array_1509_c793({a_c[715:0],793'd0},p_prime[793],c_w_793);
AND_array_1509 AND_array_1509_s793({a_s[715:0],793'd0},p_prime[793],s_w_793);
AND_array_1509 AND_array_1509_c794({a_c[714:0],794'd0},p_prime[794],c_w_794);
AND_array_1509 AND_array_1509_s794({a_s[714:0],794'd0},p_prime[794],s_w_794);
AND_array_1509 AND_array_1509_c795({a_c[713:0],795'd0},p_prime[795],c_w_795);
AND_array_1509 AND_array_1509_s795({a_s[713:0],795'd0},p_prime[795],s_w_795);
AND_array_1509 AND_array_1509_c796({a_c[712:0],796'd0},p_prime[796],c_w_796);
AND_array_1509 AND_array_1509_s796({a_s[712:0],796'd0},p_prime[796],s_w_796);
AND_array_1509 AND_array_1509_c797({a_c[711:0],797'd0},p_prime[797],c_w_797);
AND_array_1509 AND_array_1509_s797({a_s[711:0],797'd0},p_prime[797],s_w_797);
AND_array_1509 AND_array_1509_c798({a_c[710:0],798'd0},p_prime[798],c_w_798);
AND_array_1509 AND_array_1509_s798({a_s[710:0],798'd0},p_prime[798],s_w_798);
AND_array_1509 AND_array_1509_c799({a_c[709:0],799'd0},p_prime[799],c_w_799);
AND_array_1509 AND_array_1509_s799({a_s[709:0],799'd0},p_prime[799],s_w_799);
AND_array_1509 AND_array_1509_c800({a_c[708:0],800'd0},p_prime[800],c_w_800);
AND_array_1509 AND_array_1509_s800({a_s[708:0],800'd0},p_prime[800],s_w_800);
AND_array_1509 AND_array_1509_c801({a_c[707:0],801'd0},p_prime[801],c_w_801);
AND_array_1509 AND_array_1509_s801({a_s[707:0],801'd0},p_prime[801],s_w_801);
AND_array_1509 AND_array_1509_c802({a_c[706:0],802'd0},p_prime[802],c_w_802);
AND_array_1509 AND_array_1509_s802({a_s[706:0],802'd0},p_prime[802],s_w_802);
AND_array_1509 AND_array_1509_c803({a_c[705:0],803'd0},p_prime[803],c_w_803);
AND_array_1509 AND_array_1509_s803({a_s[705:0],803'd0},p_prime[803],s_w_803);
AND_array_1509 AND_array_1509_c804({a_c[704:0],804'd0},p_prime[804],c_w_804);
AND_array_1509 AND_array_1509_s804({a_s[704:0],804'd0},p_prime[804],s_w_804);
AND_array_1509 AND_array_1509_c805({a_c[703:0],805'd0},p_prime[805],c_w_805);
AND_array_1509 AND_array_1509_s805({a_s[703:0],805'd0},p_prime[805],s_w_805);
AND_array_1509 AND_array_1509_c806({a_c[702:0],806'd0},p_prime[806],c_w_806);
AND_array_1509 AND_array_1509_s806({a_s[702:0],806'd0},p_prime[806],s_w_806);
AND_array_1509 AND_array_1509_c807({a_c[701:0],807'd0},p_prime[807],c_w_807);
AND_array_1509 AND_array_1509_s807({a_s[701:0],807'd0},p_prime[807],s_w_807);
AND_array_1509 AND_array_1509_c808({a_c[700:0],808'd0},p_prime[808],c_w_808);
AND_array_1509 AND_array_1509_s808({a_s[700:0],808'd0},p_prime[808],s_w_808);
AND_array_1509 AND_array_1509_c809({a_c[699:0],809'd0},p_prime[809],c_w_809);
AND_array_1509 AND_array_1509_s809({a_s[699:0],809'd0},p_prime[809],s_w_809);
AND_array_1509 AND_array_1509_c810({a_c[698:0],810'd0},p_prime[810],c_w_810);
AND_array_1509 AND_array_1509_s810({a_s[698:0],810'd0},p_prime[810],s_w_810);
AND_array_1509 AND_array_1509_c811({a_c[697:0],811'd0},p_prime[811],c_w_811);
AND_array_1509 AND_array_1509_s811({a_s[697:0],811'd0},p_prime[811],s_w_811);
AND_array_1509 AND_array_1509_c812({a_c[696:0],812'd0},p_prime[812],c_w_812);
AND_array_1509 AND_array_1509_s812({a_s[696:0],812'd0},p_prime[812],s_w_812);
AND_array_1509 AND_array_1509_c813({a_c[695:0],813'd0},p_prime[813],c_w_813);
AND_array_1509 AND_array_1509_s813({a_s[695:0],813'd0},p_prime[813],s_w_813);
AND_array_1509 AND_array_1509_c814({a_c[694:0],814'd0},p_prime[814],c_w_814);
AND_array_1509 AND_array_1509_s814({a_s[694:0],814'd0},p_prime[814],s_w_814);
AND_array_1509 AND_array_1509_c815({a_c[693:0],815'd0},p_prime[815],c_w_815);
AND_array_1509 AND_array_1509_s815({a_s[693:0],815'd0},p_prime[815],s_w_815);
AND_array_1509 AND_array_1509_c816({a_c[692:0],816'd0},p_prime[816],c_w_816);
AND_array_1509 AND_array_1509_s816({a_s[692:0],816'd0},p_prime[816],s_w_816);
AND_array_1509 AND_array_1509_c817({a_c[691:0],817'd0},p_prime[817],c_w_817);
AND_array_1509 AND_array_1509_s817({a_s[691:0],817'd0},p_prime[817],s_w_817);
AND_array_1509 AND_array_1509_c818({a_c[690:0],818'd0},p_prime[818],c_w_818);
AND_array_1509 AND_array_1509_s818({a_s[690:0],818'd0},p_prime[818],s_w_818);
AND_array_1509 AND_array_1509_c819({a_c[689:0],819'd0},p_prime[819],c_w_819);
AND_array_1509 AND_array_1509_s819({a_s[689:0],819'd0},p_prime[819],s_w_819);
AND_array_1509 AND_array_1509_c820({a_c[688:0],820'd0},p_prime[820],c_w_820);
AND_array_1509 AND_array_1509_s820({a_s[688:0],820'd0},p_prime[820],s_w_820);
AND_array_1509 AND_array_1509_c821({a_c[687:0],821'd0},p_prime[821],c_w_821);
AND_array_1509 AND_array_1509_s821({a_s[687:0],821'd0},p_prime[821],s_w_821);
AND_array_1509 AND_array_1509_c822({a_c[686:0],822'd0},p_prime[822],c_w_822);
AND_array_1509 AND_array_1509_s822({a_s[686:0],822'd0},p_prime[822],s_w_822);
AND_array_1509 AND_array_1509_c823({a_c[685:0],823'd0},p_prime[823],c_w_823);
AND_array_1509 AND_array_1509_s823({a_s[685:0],823'd0},p_prime[823],s_w_823);
AND_array_1509 AND_array_1509_c824({a_c[684:0],824'd0},p_prime[824],c_w_824);
AND_array_1509 AND_array_1509_s824({a_s[684:0],824'd0},p_prime[824],s_w_824);
AND_array_1509 AND_array_1509_c825({a_c[683:0],825'd0},p_prime[825],c_w_825);
AND_array_1509 AND_array_1509_s825({a_s[683:0],825'd0},p_prime[825],s_w_825);
AND_array_1509 AND_array_1509_c826({a_c[682:0],826'd0},p_prime[826],c_w_826);
AND_array_1509 AND_array_1509_s826({a_s[682:0],826'd0},p_prime[826],s_w_826);
AND_array_1509 AND_array_1509_c827({a_c[681:0],827'd0},p_prime[827],c_w_827);
AND_array_1509 AND_array_1509_s827({a_s[681:0],827'd0},p_prime[827],s_w_827);
AND_array_1509 AND_array_1509_c828({a_c[680:0],828'd0},p_prime[828],c_w_828);
AND_array_1509 AND_array_1509_s828({a_s[680:0],828'd0},p_prime[828],s_w_828);
AND_array_1509 AND_array_1509_c829({a_c[679:0],829'd0},p_prime[829],c_w_829);
AND_array_1509 AND_array_1509_s829({a_s[679:0],829'd0},p_prime[829],s_w_829);
AND_array_1509 AND_array_1509_c830({a_c[678:0],830'd0},p_prime[830],c_w_830);
AND_array_1509 AND_array_1509_s830({a_s[678:0],830'd0},p_prime[830],s_w_830);
AND_array_1509 AND_array_1509_c831({a_c[677:0],831'd0},p_prime[831],c_w_831);
AND_array_1509 AND_array_1509_s831({a_s[677:0],831'd0},p_prime[831],s_w_831);
AND_array_1509 AND_array_1509_c832({a_c[676:0],832'd0},p_prime[832],c_w_832);
AND_array_1509 AND_array_1509_s832({a_s[676:0],832'd0},p_prime[832],s_w_832);
AND_array_1509 AND_array_1509_c833({a_c[675:0],833'd0},p_prime[833],c_w_833);
AND_array_1509 AND_array_1509_s833({a_s[675:0],833'd0},p_prime[833],s_w_833);
AND_array_1509 AND_array_1509_c834({a_c[674:0],834'd0},p_prime[834],c_w_834);
AND_array_1509 AND_array_1509_s834({a_s[674:0],834'd0},p_prime[834],s_w_834);
AND_array_1509 AND_array_1509_c835({a_c[673:0],835'd0},p_prime[835],c_w_835);
AND_array_1509 AND_array_1509_s835({a_s[673:0],835'd0},p_prime[835],s_w_835);
AND_array_1509 AND_array_1509_c836({a_c[672:0],836'd0},p_prime[836],c_w_836);
AND_array_1509 AND_array_1509_s836({a_s[672:0],836'd0},p_prime[836],s_w_836);
AND_array_1509 AND_array_1509_c837({a_c[671:0],837'd0},p_prime[837],c_w_837);
AND_array_1509 AND_array_1509_s837({a_s[671:0],837'd0},p_prime[837],s_w_837);
AND_array_1509 AND_array_1509_c838({a_c[670:0],838'd0},p_prime[838],c_w_838);
AND_array_1509 AND_array_1509_s838({a_s[670:0],838'd0},p_prime[838],s_w_838);
AND_array_1509 AND_array_1509_c839({a_c[669:0],839'd0},p_prime[839],c_w_839);
AND_array_1509 AND_array_1509_s839({a_s[669:0],839'd0},p_prime[839],s_w_839);
AND_array_1509 AND_array_1509_c840({a_c[668:0],840'd0},p_prime[840],c_w_840);
AND_array_1509 AND_array_1509_s840({a_s[668:0],840'd0},p_prime[840],s_w_840);
AND_array_1509 AND_array_1509_c841({a_c[667:0],841'd0},p_prime[841],c_w_841);
AND_array_1509 AND_array_1509_s841({a_s[667:0],841'd0},p_prime[841],s_w_841);
AND_array_1509 AND_array_1509_c842({a_c[666:0],842'd0},p_prime[842],c_w_842);
AND_array_1509 AND_array_1509_s842({a_s[666:0],842'd0},p_prime[842],s_w_842);
AND_array_1509 AND_array_1509_c843({a_c[665:0],843'd0},p_prime[843],c_w_843);
AND_array_1509 AND_array_1509_s843({a_s[665:0],843'd0},p_prime[843],s_w_843);
AND_array_1509 AND_array_1509_c844({a_c[664:0],844'd0},p_prime[844],c_w_844);
AND_array_1509 AND_array_1509_s844({a_s[664:0],844'd0},p_prime[844],s_w_844);
AND_array_1509 AND_array_1509_c845({a_c[663:0],845'd0},p_prime[845],c_w_845);
AND_array_1509 AND_array_1509_s845({a_s[663:0],845'd0},p_prime[845],s_w_845);
AND_array_1509 AND_array_1509_c846({a_c[662:0],846'd0},p_prime[846],c_w_846);
AND_array_1509 AND_array_1509_s846({a_s[662:0],846'd0},p_prime[846],s_w_846);
AND_array_1509 AND_array_1509_c847({a_c[661:0],847'd0},p_prime[847],c_w_847);
AND_array_1509 AND_array_1509_s847({a_s[661:0],847'd0},p_prime[847],s_w_847);
AND_array_1509 AND_array_1509_c848({a_c[660:0],848'd0},p_prime[848],c_w_848);
AND_array_1509 AND_array_1509_s848({a_s[660:0],848'd0},p_prime[848],s_w_848);
AND_array_1509 AND_array_1509_c849({a_c[659:0],849'd0},p_prime[849],c_w_849);
AND_array_1509 AND_array_1509_s849({a_s[659:0],849'd0},p_prime[849],s_w_849);
AND_array_1509 AND_array_1509_c850({a_c[658:0],850'd0},p_prime[850],c_w_850);
AND_array_1509 AND_array_1509_s850({a_s[658:0],850'd0},p_prime[850],s_w_850);
AND_array_1509 AND_array_1509_c851({a_c[657:0],851'd0},p_prime[851],c_w_851);
AND_array_1509 AND_array_1509_s851({a_s[657:0],851'd0},p_prime[851],s_w_851);
AND_array_1509 AND_array_1509_c852({a_c[656:0],852'd0},p_prime[852],c_w_852);
AND_array_1509 AND_array_1509_s852({a_s[656:0],852'd0},p_prime[852],s_w_852);
AND_array_1509 AND_array_1509_c853({a_c[655:0],853'd0},p_prime[853],c_w_853);
AND_array_1509 AND_array_1509_s853({a_s[655:0],853'd0},p_prime[853],s_w_853);
AND_array_1509 AND_array_1509_c854({a_c[654:0],854'd0},p_prime[854],c_w_854);
AND_array_1509 AND_array_1509_s854({a_s[654:0],854'd0},p_prime[854],s_w_854);
AND_array_1509 AND_array_1509_c855({a_c[653:0],855'd0},p_prime[855],c_w_855);
AND_array_1509 AND_array_1509_s855({a_s[653:0],855'd0},p_prime[855],s_w_855);
AND_array_1509 AND_array_1509_c856({a_c[652:0],856'd0},p_prime[856],c_w_856);
AND_array_1509 AND_array_1509_s856({a_s[652:0],856'd0},p_prime[856],s_w_856);
AND_array_1509 AND_array_1509_c857({a_c[651:0],857'd0},p_prime[857],c_w_857);
AND_array_1509 AND_array_1509_s857({a_s[651:0],857'd0},p_prime[857],s_w_857);
AND_array_1509 AND_array_1509_c858({a_c[650:0],858'd0},p_prime[858],c_w_858);
AND_array_1509 AND_array_1509_s858({a_s[650:0],858'd0},p_prime[858],s_w_858);
AND_array_1509 AND_array_1509_c859({a_c[649:0],859'd0},p_prime[859],c_w_859);
AND_array_1509 AND_array_1509_s859({a_s[649:0],859'd0},p_prime[859],s_w_859);
AND_array_1509 AND_array_1509_c860({a_c[648:0],860'd0},p_prime[860],c_w_860);
AND_array_1509 AND_array_1509_s860({a_s[648:0],860'd0},p_prime[860],s_w_860);
AND_array_1509 AND_array_1509_c861({a_c[647:0],861'd0},p_prime[861],c_w_861);
AND_array_1509 AND_array_1509_s861({a_s[647:0],861'd0},p_prime[861],s_w_861);
AND_array_1509 AND_array_1509_c862({a_c[646:0],862'd0},p_prime[862],c_w_862);
AND_array_1509 AND_array_1509_s862({a_s[646:0],862'd0},p_prime[862],s_w_862);
AND_array_1509 AND_array_1509_c863({a_c[645:0],863'd0},p_prime[863],c_w_863);
AND_array_1509 AND_array_1509_s863({a_s[645:0],863'd0},p_prime[863],s_w_863);
AND_array_1509 AND_array_1509_c864({a_c[644:0],864'd0},p_prime[864],c_w_864);
AND_array_1509 AND_array_1509_s864({a_s[644:0],864'd0},p_prime[864],s_w_864);
AND_array_1509 AND_array_1509_c865({a_c[643:0],865'd0},p_prime[865],c_w_865);
AND_array_1509 AND_array_1509_s865({a_s[643:0],865'd0},p_prime[865],s_w_865);
AND_array_1509 AND_array_1509_c866({a_c[642:0],866'd0},p_prime[866],c_w_866);
AND_array_1509 AND_array_1509_s866({a_s[642:0],866'd0},p_prime[866],s_w_866);
AND_array_1509 AND_array_1509_c867({a_c[641:0],867'd0},p_prime[867],c_w_867);
AND_array_1509 AND_array_1509_s867({a_s[641:0],867'd0},p_prime[867],s_w_867);
AND_array_1509 AND_array_1509_c868({a_c[640:0],868'd0},p_prime[868],c_w_868);
AND_array_1509 AND_array_1509_s868({a_s[640:0],868'd0},p_prime[868],s_w_868);
AND_array_1509 AND_array_1509_c869({a_c[639:0],869'd0},p_prime[869],c_w_869);
AND_array_1509 AND_array_1509_s869({a_s[639:0],869'd0},p_prime[869],s_w_869);
AND_array_1509 AND_array_1509_c870({a_c[638:0],870'd0},p_prime[870],c_w_870);
AND_array_1509 AND_array_1509_s870({a_s[638:0],870'd0},p_prime[870],s_w_870);
AND_array_1509 AND_array_1509_c871({a_c[637:0],871'd0},p_prime[871],c_w_871);
AND_array_1509 AND_array_1509_s871({a_s[637:0],871'd0},p_prime[871],s_w_871);
AND_array_1509 AND_array_1509_c872({a_c[636:0],872'd0},p_prime[872],c_w_872);
AND_array_1509 AND_array_1509_s872({a_s[636:0],872'd0},p_prime[872],s_w_872);
AND_array_1509 AND_array_1509_c873({a_c[635:0],873'd0},p_prime[873],c_w_873);
AND_array_1509 AND_array_1509_s873({a_s[635:0],873'd0},p_prime[873],s_w_873);
AND_array_1509 AND_array_1509_c874({a_c[634:0],874'd0},p_prime[874],c_w_874);
AND_array_1509 AND_array_1509_s874({a_s[634:0],874'd0},p_prime[874],s_w_874);
AND_array_1509 AND_array_1509_c875({a_c[633:0],875'd0},p_prime[875],c_w_875);
AND_array_1509 AND_array_1509_s875({a_s[633:0],875'd0},p_prime[875],s_w_875);
AND_array_1509 AND_array_1509_c876({a_c[632:0],876'd0},p_prime[876],c_w_876);
AND_array_1509 AND_array_1509_s876({a_s[632:0],876'd0},p_prime[876],s_w_876);
AND_array_1509 AND_array_1509_c877({a_c[631:0],877'd0},p_prime[877],c_w_877);
AND_array_1509 AND_array_1509_s877({a_s[631:0],877'd0},p_prime[877],s_w_877);
AND_array_1509 AND_array_1509_c878({a_c[630:0],878'd0},p_prime[878],c_w_878);
AND_array_1509 AND_array_1509_s878({a_s[630:0],878'd0},p_prime[878],s_w_878);
AND_array_1509 AND_array_1509_c879({a_c[629:0],879'd0},p_prime[879],c_w_879);
AND_array_1509 AND_array_1509_s879({a_s[629:0],879'd0},p_prime[879],s_w_879);
AND_array_1509 AND_array_1509_c880({a_c[628:0],880'd0},p_prime[880],c_w_880);
AND_array_1509 AND_array_1509_s880({a_s[628:0],880'd0},p_prime[880],s_w_880);
AND_array_1509 AND_array_1509_c881({a_c[627:0],881'd0},p_prime[881],c_w_881);
AND_array_1509 AND_array_1509_s881({a_s[627:0],881'd0},p_prime[881],s_w_881);
AND_array_1509 AND_array_1509_c882({a_c[626:0],882'd0},p_prime[882],c_w_882);
AND_array_1509 AND_array_1509_s882({a_s[626:0],882'd0},p_prime[882],s_w_882);
AND_array_1509 AND_array_1509_c883({a_c[625:0],883'd0},p_prime[883],c_w_883);
AND_array_1509 AND_array_1509_s883({a_s[625:0],883'd0},p_prime[883],s_w_883);
AND_array_1509 AND_array_1509_c884({a_c[624:0],884'd0},p_prime[884],c_w_884);
AND_array_1509 AND_array_1509_s884({a_s[624:0],884'd0},p_prime[884],s_w_884);
AND_array_1509 AND_array_1509_c885({a_c[623:0],885'd0},p_prime[885],c_w_885);
AND_array_1509 AND_array_1509_s885({a_s[623:0],885'd0},p_prime[885],s_w_885);
AND_array_1509 AND_array_1509_c886({a_c[622:0],886'd0},p_prime[886],c_w_886);
AND_array_1509 AND_array_1509_s886({a_s[622:0],886'd0},p_prime[886],s_w_886);
AND_array_1509 AND_array_1509_c887({a_c[621:0],887'd0},p_prime[887],c_w_887);
AND_array_1509 AND_array_1509_s887({a_s[621:0],887'd0},p_prime[887],s_w_887);
AND_array_1509 AND_array_1509_c888({a_c[620:0],888'd0},p_prime[888],c_w_888);
AND_array_1509 AND_array_1509_s888({a_s[620:0],888'd0},p_prime[888],s_w_888);
AND_array_1509 AND_array_1509_c889({a_c[619:0],889'd0},p_prime[889],c_w_889);
AND_array_1509 AND_array_1509_s889({a_s[619:0],889'd0},p_prime[889],s_w_889);
AND_array_1509 AND_array_1509_c890({a_c[618:0],890'd0},p_prime[890],c_w_890);
AND_array_1509 AND_array_1509_s890({a_s[618:0],890'd0},p_prime[890],s_w_890);
AND_array_1509 AND_array_1509_c891({a_c[617:0],891'd0},p_prime[891],c_w_891);
AND_array_1509 AND_array_1509_s891({a_s[617:0],891'd0},p_prime[891],s_w_891);
AND_array_1509 AND_array_1509_c892({a_c[616:0],892'd0},p_prime[892],c_w_892);
AND_array_1509 AND_array_1509_s892({a_s[616:0],892'd0},p_prime[892],s_w_892);
AND_array_1509 AND_array_1509_c893({a_c[615:0],893'd0},p_prime[893],c_w_893);
AND_array_1509 AND_array_1509_s893({a_s[615:0],893'd0},p_prime[893],s_w_893);
AND_array_1509 AND_array_1509_c894({a_c[614:0],894'd0},p_prime[894],c_w_894);
AND_array_1509 AND_array_1509_s894({a_s[614:0],894'd0},p_prime[894],s_w_894);
AND_array_1509 AND_array_1509_c895({a_c[613:0],895'd0},p_prime[895],c_w_895);
AND_array_1509 AND_array_1509_s895({a_s[613:0],895'd0},p_prime[895],s_w_895);
AND_array_1509 AND_array_1509_c896({a_c[612:0],896'd0},p_prime[896],c_w_896);
AND_array_1509 AND_array_1509_s896({a_s[612:0],896'd0},p_prime[896],s_w_896);
AND_array_1509 AND_array_1509_c897({a_c[611:0],897'd0},p_prime[897],c_w_897);
AND_array_1509 AND_array_1509_s897({a_s[611:0],897'd0},p_prime[897],s_w_897);
AND_array_1509 AND_array_1509_c898({a_c[610:0],898'd0},p_prime[898],c_w_898);
AND_array_1509 AND_array_1509_s898({a_s[610:0],898'd0},p_prime[898],s_w_898);
AND_array_1509 AND_array_1509_c899({a_c[609:0],899'd0},p_prime[899],c_w_899);
AND_array_1509 AND_array_1509_s899({a_s[609:0],899'd0},p_prime[899],s_w_899);
AND_array_1509 AND_array_1509_c900({a_c[608:0],900'd0},p_prime[900],c_w_900);
AND_array_1509 AND_array_1509_s900({a_s[608:0],900'd0},p_prime[900],s_w_900);
AND_array_1509 AND_array_1509_c901({a_c[607:0],901'd0},p_prime[901],c_w_901);
AND_array_1509 AND_array_1509_s901({a_s[607:0],901'd0},p_prime[901],s_w_901);
AND_array_1509 AND_array_1509_c902({a_c[606:0],902'd0},p_prime[902],c_w_902);
AND_array_1509 AND_array_1509_s902({a_s[606:0],902'd0},p_prime[902],s_w_902);
AND_array_1509 AND_array_1509_c903({a_c[605:0],903'd0},p_prime[903],c_w_903);
AND_array_1509 AND_array_1509_s903({a_s[605:0],903'd0},p_prime[903],s_w_903);
AND_array_1509 AND_array_1509_c904({a_c[604:0],904'd0},p_prime[904],c_w_904);
AND_array_1509 AND_array_1509_s904({a_s[604:0],904'd0},p_prime[904],s_w_904);
AND_array_1509 AND_array_1509_c905({a_c[603:0],905'd0},p_prime[905],c_w_905);
AND_array_1509 AND_array_1509_s905({a_s[603:0],905'd0},p_prime[905],s_w_905);
AND_array_1509 AND_array_1509_c906({a_c[602:0],906'd0},p_prime[906],c_w_906);
AND_array_1509 AND_array_1509_s906({a_s[602:0],906'd0},p_prime[906],s_w_906);
AND_array_1509 AND_array_1509_c907({a_c[601:0],907'd0},p_prime[907],c_w_907);
AND_array_1509 AND_array_1509_s907({a_s[601:0],907'd0},p_prime[907],s_w_907);
AND_array_1509 AND_array_1509_c908({a_c[600:0],908'd0},p_prime[908],c_w_908);
AND_array_1509 AND_array_1509_s908({a_s[600:0],908'd0},p_prime[908],s_w_908);
AND_array_1509 AND_array_1509_c909({a_c[599:0],909'd0},p_prime[909],c_w_909);
AND_array_1509 AND_array_1509_s909({a_s[599:0],909'd0},p_prime[909],s_w_909);
AND_array_1509 AND_array_1509_c910({a_c[598:0],910'd0},p_prime[910],c_w_910);
AND_array_1509 AND_array_1509_s910({a_s[598:0],910'd0},p_prime[910],s_w_910);
AND_array_1509 AND_array_1509_c911({a_c[597:0],911'd0},p_prime[911],c_w_911);
AND_array_1509 AND_array_1509_s911({a_s[597:0],911'd0},p_prime[911],s_w_911);
AND_array_1509 AND_array_1509_c912({a_c[596:0],912'd0},p_prime[912],c_w_912);
AND_array_1509 AND_array_1509_s912({a_s[596:0],912'd0},p_prime[912],s_w_912);
AND_array_1509 AND_array_1509_c913({a_c[595:0],913'd0},p_prime[913],c_w_913);
AND_array_1509 AND_array_1509_s913({a_s[595:0],913'd0},p_prime[913],s_w_913);
AND_array_1509 AND_array_1509_c914({a_c[594:0],914'd0},p_prime[914],c_w_914);
AND_array_1509 AND_array_1509_s914({a_s[594:0],914'd0},p_prime[914],s_w_914);
AND_array_1509 AND_array_1509_c915({a_c[593:0],915'd0},p_prime[915],c_w_915);
AND_array_1509 AND_array_1509_s915({a_s[593:0],915'd0},p_prime[915],s_w_915);
AND_array_1509 AND_array_1509_c916({a_c[592:0],916'd0},p_prime[916],c_w_916);
AND_array_1509 AND_array_1509_s916({a_s[592:0],916'd0},p_prime[916],s_w_916);
AND_array_1509 AND_array_1509_c917({a_c[591:0],917'd0},p_prime[917],c_w_917);
AND_array_1509 AND_array_1509_s917({a_s[591:0],917'd0},p_prime[917],s_w_917);
AND_array_1509 AND_array_1509_c918({a_c[590:0],918'd0},p_prime[918],c_w_918);
AND_array_1509 AND_array_1509_s918({a_s[590:0],918'd0},p_prime[918],s_w_918);
AND_array_1509 AND_array_1509_c919({a_c[589:0],919'd0},p_prime[919],c_w_919);
AND_array_1509 AND_array_1509_s919({a_s[589:0],919'd0},p_prime[919],s_w_919);
AND_array_1509 AND_array_1509_c920({a_c[588:0],920'd0},p_prime[920],c_w_920);
AND_array_1509 AND_array_1509_s920({a_s[588:0],920'd0},p_prime[920],s_w_920);
AND_array_1509 AND_array_1509_c921({a_c[587:0],921'd0},p_prime[921],c_w_921);
AND_array_1509 AND_array_1509_s921({a_s[587:0],921'd0},p_prime[921],s_w_921);
AND_array_1509 AND_array_1509_c922({a_c[586:0],922'd0},p_prime[922],c_w_922);
AND_array_1509 AND_array_1509_s922({a_s[586:0],922'd0},p_prime[922],s_w_922);
AND_array_1509 AND_array_1509_c923({a_c[585:0],923'd0},p_prime[923],c_w_923);
AND_array_1509 AND_array_1509_s923({a_s[585:0],923'd0},p_prime[923],s_w_923);
AND_array_1509 AND_array_1509_c924({a_c[584:0],924'd0},p_prime[924],c_w_924);
AND_array_1509 AND_array_1509_s924({a_s[584:0],924'd0},p_prime[924],s_w_924);
AND_array_1509 AND_array_1509_c925({a_c[583:0],925'd0},p_prime[925],c_w_925);
AND_array_1509 AND_array_1509_s925({a_s[583:0],925'd0},p_prime[925],s_w_925);
AND_array_1509 AND_array_1509_c926({a_c[582:0],926'd0},p_prime[926],c_w_926);
AND_array_1509 AND_array_1509_s926({a_s[582:0],926'd0},p_prime[926],s_w_926);
AND_array_1509 AND_array_1509_c927({a_c[581:0],927'd0},p_prime[927],c_w_927);
AND_array_1509 AND_array_1509_s927({a_s[581:0],927'd0},p_prime[927],s_w_927);
AND_array_1509 AND_array_1509_c928({a_c[580:0],928'd0},p_prime[928],c_w_928);
AND_array_1509 AND_array_1509_s928({a_s[580:0],928'd0},p_prime[928],s_w_928);
AND_array_1509 AND_array_1509_c929({a_c[579:0],929'd0},p_prime[929],c_w_929);
AND_array_1509 AND_array_1509_s929({a_s[579:0],929'd0},p_prime[929],s_w_929);
AND_array_1509 AND_array_1509_c930({a_c[578:0],930'd0},p_prime[930],c_w_930);
AND_array_1509 AND_array_1509_s930({a_s[578:0],930'd0},p_prime[930],s_w_930);
AND_array_1509 AND_array_1509_c931({a_c[577:0],931'd0},p_prime[931],c_w_931);
AND_array_1509 AND_array_1509_s931({a_s[577:0],931'd0},p_prime[931],s_w_931);
AND_array_1509 AND_array_1509_c932({a_c[576:0],932'd0},p_prime[932],c_w_932);
AND_array_1509 AND_array_1509_s932({a_s[576:0],932'd0},p_prime[932],s_w_932);
AND_array_1509 AND_array_1509_c933({a_c[575:0],933'd0},p_prime[933],c_w_933);
AND_array_1509 AND_array_1509_s933({a_s[575:0],933'd0},p_prime[933],s_w_933);
AND_array_1509 AND_array_1509_c934({a_c[574:0],934'd0},p_prime[934],c_w_934);
AND_array_1509 AND_array_1509_s934({a_s[574:0],934'd0},p_prime[934],s_w_934);
AND_array_1509 AND_array_1509_c935({a_c[573:0],935'd0},p_prime[935],c_w_935);
AND_array_1509 AND_array_1509_s935({a_s[573:0],935'd0},p_prime[935],s_w_935);
AND_array_1509 AND_array_1509_c936({a_c[572:0],936'd0},p_prime[936],c_w_936);
AND_array_1509 AND_array_1509_s936({a_s[572:0],936'd0},p_prime[936],s_w_936);
AND_array_1509 AND_array_1509_c937({a_c[571:0],937'd0},p_prime[937],c_w_937);
AND_array_1509 AND_array_1509_s937({a_s[571:0],937'd0},p_prime[937],s_w_937);
AND_array_1509 AND_array_1509_c938({a_c[570:0],938'd0},p_prime[938],c_w_938);
AND_array_1509 AND_array_1509_s938({a_s[570:0],938'd0},p_prime[938],s_w_938);
AND_array_1509 AND_array_1509_c939({a_c[569:0],939'd0},p_prime[939],c_w_939);
AND_array_1509 AND_array_1509_s939({a_s[569:0],939'd0},p_prime[939],s_w_939);
AND_array_1509 AND_array_1509_c940({a_c[568:0],940'd0},p_prime[940],c_w_940);
AND_array_1509 AND_array_1509_s940({a_s[568:0],940'd0},p_prime[940],s_w_940);
AND_array_1509 AND_array_1509_c941({a_c[567:0],941'd0},p_prime[941],c_w_941);
AND_array_1509 AND_array_1509_s941({a_s[567:0],941'd0},p_prime[941],s_w_941);
AND_array_1509 AND_array_1509_c942({a_c[566:0],942'd0},p_prime[942],c_w_942);
AND_array_1509 AND_array_1509_s942({a_s[566:0],942'd0},p_prime[942],s_w_942);
AND_array_1509 AND_array_1509_c943({a_c[565:0],943'd0},p_prime[943],c_w_943);
AND_array_1509 AND_array_1509_s943({a_s[565:0],943'd0},p_prime[943],s_w_943);
AND_array_1509 AND_array_1509_c944({a_c[564:0],944'd0},p_prime[944],c_w_944);
AND_array_1509 AND_array_1509_s944({a_s[564:0],944'd0},p_prime[944],s_w_944);
AND_array_1509 AND_array_1509_c945({a_c[563:0],945'd0},p_prime[945],c_w_945);
AND_array_1509 AND_array_1509_s945({a_s[563:0],945'd0},p_prime[945],s_w_945);
AND_array_1509 AND_array_1509_c946({a_c[562:0],946'd0},p_prime[946],c_w_946);
AND_array_1509 AND_array_1509_s946({a_s[562:0],946'd0},p_prime[946],s_w_946);
AND_array_1509 AND_array_1509_c947({a_c[561:0],947'd0},p_prime[947],c_w_947);
AND_array_1509 AND_array_1509_s947({a_s[561:0],947'd0},p_prime[947],s_w_947);
AND_array_1509 AND_array_1509_c948({a_c[560:0],948'd0},p_prime[948],c_w_948);
AND_array_1509 AND_array_1509_s948({a_s[560:0],948'd0},p_prime[948],s_w_948);
AND_array_1509 AND_array_1509_c949({a_c[559:0],949'd0},p_prime[949],c_w_949);
AND_array_1509 AND_array_1509_s949({a_s[559:0],949'd0},p_prime[949],s_w_949);
AND_array_1509 AND_array_1509_c950({a_c[558:0],950'd0},p_prime[950],c_w_950);
AND_array_1509 AND_array_1509_s950({a_s[558:0],950'd0},p_prime[950],s_w_950);
AND_array_1509 AND_array_1509_c951({a_c[557:0],951'd0},p_prime[951],c_w_951);
AND_array_1509 AND_array_1509_s951({a_s[557:0],951'd0},p_prime[951],s_w_951);
AND_array_1509 AND_array_1509_c952({a_c[556:0],952'd0},p_prime[952],c_w_952);
AND_array_1509 AND_array_1509_s952({a_s[556:0],952'd0},p_prime[952],s_w_952);
AND_array_1509 AND_array_1509_c953({a_c[555:0],953'd0},p_prime[953],c_w_953);
AND_array_1509 AND_array_1509_s953({a_s[555:0],953'd0},p_prime[953],s_w_953);
AND_array_1509 AND_array_1509_c954({a_c[554:0],954'd0},p_prime[954],c_w_954);
AND_array_1509 AND_array_1509_s954({a_s[554:0],954'd0},p_prime[954],s_w_954);
AND_array_1509 AND_array_1509_c955({a_c[553:0],955'd0},p_prime[955],c_w_955);
AND_array_1509 AND_array_1509_s955({a_s[553:0],955'd0},p_prime[955],s_w_955);
AND_array_1509 AND_array_1509_c956({a_c[552:0],956'd0},p_prime[956],c_w_956);
AND_array_1509 AND_array_1509_s956({a_s[552:0],956'd0},p_prime[956],s_w_956);
AND_array_1509 AND_array_1509_c957({a_c[551:0],957'd0},p_prime[957],c_w_957);
AND_array_1509 AND_array_1509_s957({a_s[551:0],957'd0},p_prime[957],s_w_957);
AND_array_1509 AND_array_1509_c958({a_c[550:0],958'd0},p_prime[958],c_w_958);
AND_array_1509 AND_array_1509_s958({a_s[550:0],958'd0},p_prime[958],s_w_958);
AND_array_1509 AND_array_1509_c959({a_c[549:0],959'd0},p_prime[959],c_w_959);
AND_array_1509 AND_array_1509_s959({a_s[549:0],959'd0},p_prime[959],s_w_959);
AND_array_1509 AND_array_1509_c960({a_c[548:0],960'd0},p_prime[960],c_w_960);
AND_array_1509 AND_array_1509_s960({a_s[548:0],960'd0},p_prime[960],s_w_960);
AND_array_1509 AND_array_1509_c961({a_c[547:0],961'd0},p_prime[961],c_w_961);
AND_array_1509 AND_array_1509_s961({a_s[547:0],961'd0},p_prime[961],s_w_961);
AND_array_1509 AND_array_1509_c962({a_c[546:0],962'd0},p_prime[962],c_w_962);
AND_array_1509 AND_array_1509_s962({a_s[546:0],962'd0},p_prime[962],s_w_962);
AND_array_1509 AND_array_1509_c963({a_c[545:0],963'd0},p_prime[963],c_w_963);
AND_array_1509 AND_array_1509_s963({a_s[545:0],963'd0},p_prime[963],s_w_963);
AND_array_1509 AND_array_1509_c964({a_c[544:0],964'd0},p_prime[964],c_w_964);
AND_array_1509 AND_array_1509_s964({a_s[544:0],964'd0},p_prime[964],s_w_964);
AND_array_1509 AND_array_1509_c965({a_c[543:0],965'd0},p_prime[965],c_w_965);
AND_array_1509 AND_array_1509_s965({a_s[543:0],965'd0},p_prime[965],s_w_965);
AND_array_1509 AND_array_1509_c966({a_c[542:0],966'd0},p_prime[966],c_w_966);
AND_array_1509 AND_array_1509_s966({a_s[542:0],966'd0},p_prime[966],s_w_966);
AND_array_1509 AND_array_1509_c967({a_c[541:0],967'd0},p_prime[967],c_w_967);
AND_array_1509 AND_array_1509_s967({a_s[541:0],967'd0},p_prime[967],s_w_967);
AND_array_1509 AND_array_1509_c968({a_c[540:0],968'd0},p_prime[968],c_w_968);
AND_array_1509 AND_array_1509_s968({a_s[540:0],968'd0},p_prime[968],s_w_968);
AND_array_1509 AND_array_1509_c969({a_c[539:0],969'd0},p_prime[969],c_w_969);
AND_array_1509 AND_array_1509_s969({a_s[539:0],969'd0},p_prime[969],s_w_969);
AND_array_1509 AND_array_1509_c970({a_c[538:0],970'd0},p_prime[970],c_w_970);
AND_array_1509 AND_array_1509_s970({a_s[538:0],970'd0},p_prime[970],s_w_970);
AND_array_1509 AND_array_1509_c971({a_c[537:0],971'd0},p_prime[971],c_w_971);
AND_array_1509 AND_array_1509_s971({a_s[537:0],971'd0},p_prime[971],s_w_971);
AND_array_1509 AND_array_1509_c972({a_c[536:0],972'd0},p_prime[972],c_w_972);
AND_array_1509 AND_array_1509_s972({a_s[536:0],972'd0},p_prime[972],s_w_972);
AND_array_1509 AND_array_1509_c973({a_c[535:0],973'd0},p_prime[973],c_w_973);
AND_array_1509 AND_array_1509_s973({a_s[535:0],973'd0},p_prime[973],s_w_973);
AND_array_1509 AND_array_1509_c974({a_c[534:0],974'd0},p_prime[974],c_w_974);
AND_array_1509 AND_array_1509_s974({a_s[534:0],974'd0},p_prime[974],s_w_974);
AND_array_1509 AND_array_1509_c975({a_c[533:0],975'd0},p_prime[975],c_w_975);
AND_array_1509 AND_array_1509_s975({a_s[533:0],975'd0},p_prime[975],s_w_975);
AND_array_1509 AND_array_1509_c976({a_c[532:0],976'd0},p_prime[976],c_w_976);
AND_array_1509 AND_array_1509_s976({a_s[532:0],976'd0},p_prime[976],s_w_976);
AND_array_1509 AND_array_1509_c977({a_c[531:0],977'd0},p_prime[977],c_w_977);
AND_array_1509 AND_array_1509_s977({a_s[531:0],977'd0},p_prime[977],s_w_977);
AND_array_1509 AND_array_1509_c978({a_c[530:0],978'd0},p_prime[978],c_w_978);
AND_array_1509 AND_array_1509_s978({a_s[530:0],978'd0},p_prime[978],s_w_978);
AND_array_1509 AND_array_1509_c979({a_c[529:0],979'd0},p_prime[979],c_w_979);
AND_array_1509 AND_array_1509_s979({a_s[529:0],979'd0},p_prime[979],s_w_979);
AND_array_1509 AND_array_1509_c980({a_c[528:0],980'd0},p_prime[980],c_w_980);
AND_array_1509 AND_array_1509_s980({a_s[528:0],980'd0},p_prime[980],s_w_980);
AND_array_1509 AND_array_1509_c981({a_c[527:0],981'd0},p_prime[981],c_w_981);
AND_array_1509 AND_array_1509_s981({a_s[527:0],981'd0},p_prime[981],s_w_981);
AND_array_1509 AND_array_1509_c982({a_c[526:0],982'd0},p_prime[982],c_w_982);
AND_array_1509 AND_array_1509_s982({a_s[526:0],982'd0},p_prime[982],s_w_982);
AND_array_1509 AND_array_1509_c983({a_c[525:0],983'd0},p_prime[983],c_w_983);
AND_array_1509 AND_array_1509_s983({a_s[525:0],983'd0},p_prime[983],s_w_983);
AND_array_1509 AND_array_1509_c984({a_c[524:0],984'd0},p_prime[984],c_w_984);
AND_array_1509 AND_array_1509_s984({a_s[524:0],984'd0},p_prime[984],s_w_984);
AND_array_1509 AND_array_1509_c985({a_c[523:0],985'd0},p_prime[985],c_w_985);
AND_array_1509 AND_array_1509_s985({a_s[523:0],985'd0},p_prime[985],s_w_985);
AND_array_1509 AND_array_1509_c986({a_c[522:0],986'd0},p_prime[986],c_w_986);
AND_array_1509 AND_array_1509_s986({a_s[522:0],986'd0},p_prime[986],s_w_986);
AND_array_1509 AND_array_1509_c987({a_c[521:0],987'd0},p_prime[987],c_w_987);
AND_array_1509 AND_array_1509_s987({a_s[521:0],987'd0},p_prime[987],s_w_987);
AND_array_1509 AND_array_1509_c988({a_c[520:0],988'd0},p_prime[988],c_w_988);
AND_array_1509 AND_array_1509_s988({a_s[520:0],988'd0},p_prime[988],s_w_988);
AND_array_1509 AND_array_1509_c989({a_c[519:0],989'd0},p_prime[989],c_w_989);
AND_array_1509 AND_array_1509_s989({a_s[519:0],989'd0},p_prime[989],s_w_989);
AND_array_1509 AND_array_1509_c990({a_c[518:0],990'd0},p_prime[990],c_w_990);
AND_array_1509 AND_array_1509_s990({a_s[518:0],990'd0},p_prime[990],s_w_990);
AND_array_1509 AND_array_1509_c991({a_c[517:0],991'd0},p_prime[991],c_w_991);
AND_array_1509 AND_array_1509_s991({a_s[517:0],991'd0},p_prime[991],s_w_991);
AND_array_1509 AND_array_1509_c992({a_c[516:0],992'd0},p_prime[992],c_w_992);
AND_array_1509 AND_array_1509_s992({a_s[516:0],992'd0},p_prime[992],s_w_992);
AND_array_1509 AND_array_1509_c993({a_c[515:0],993'd0},p_prime[993],c_w_993);
AND_array_1509 AND_array_1509_s993({a_s[515:0],993'd0},p_prime[993],s_w_993);
AND_array_1509 AND_array_1509_c994({a_c[514:0],994'd0},p_prime[994],c_w_994);
AND_array_1509 AND_array_1509_s994({a_s[514:0],994'd0},p_prime[994],s_w_994);
AND_array_1509 AND_array_1509_c995({a_c[513:0],995'd0},p_prime[995],c_w_995);
AND_array_1509 AND_array_1509_s995({a_s[513:0],995'd0},p_prime[995],s_w_995);
AND_array_1509 AND_array_1509_c996({a_c[512:0],996'd0},p_prime[996],c_w_996);
AND_array_1509 AND_array_1509_s996({a_s[512:0],996'd0},p_prime[996],s_w_996);
AND_array_1509 AND_array_1509_c997({a_c[511:0],997'd0},p_prime[997],c_w_997);
AND_array_1509 AND_array_1509_s997({a_s[511:0],997'd0},p_prime[997],s_w_997);
AND_array_1509 AND_array_1509_c998({a_c[510:0],998'd0},p_prime[998],c_w_998);
AND_array_1509 AND_array_1509_s998({a_s[510:0],998'd0},p_prime[998],s_w_998);
AND_array_1509 AND_array_1509_c999({a_c[509:0],999'd0},p_prime[999],c_w_999);
AND_array_1509 AND_array_1509_s999({a_s[509:0],999'd0},p_prime[999],s_w_999);
AND_array_1509 AND_array_1509_c1000({a_c[508:0],1000'd0},p_prime[1000],c_w_1000);
AND_array_1509 AND_array_1509_s1000({a_s[508:0],1000'd0},p_prime[1000],s_w_1000);
AND_array_1509 AND_array_1509_c1001({a_c[507:0],1001'd0},p_prime[1001],c_w_1001);
AND_array_1509 AND_array_1509_s1001({a_s[507:0],1001'd0},p_prime[1001],s_w_1001);
AND_array_1509 AND_array_1509_c1002({a_c[506:0],1002'd0},p_prime[1002],c_w_1002);
AND_array_1509 AND_array_1509_s1002({a_s[506:0],1002'd0},p_prime[1002],s_w_1002);
AND_array_1509 AND_array_1509_c1003({a_c[505:0],1003'd0},p_prime[1003],c_w_1003);
AND_array_1509 AND_array_1509_s1003({a_s[505:0],1003'd0},p_prime[1003],s_w_1003);
AND_array_1509 AND_array_1509_c1004({a_c[504:0],1004'd0},p_prime[1004],c_w_1004);
AND_array_1509 AND_array_1509_s1004({a_s[504:0],1004'd0},p_prime[1004],s_w_1004);
AND_array_1509 AND_array_1509_c1005({a_c[503:0],1005'd0},p_prime[1005],c_w_1005);
AND_array_1509 AND_array_1509_s1005({a_s[503:0],1005'd0},p_prime[1005],s_w_1005);
AND_array_1509 AND_array_1509_c1006({a_c[502:0],1006'd0},p_prime[1006],c_w_1006);
AND_array_1509 AND_array_1509_s1006({a_s[502:0],1006'd0},p_prime[1006],s_w_1006);
AND_array_1509 AND_array_1509_c1007({a_c[501:0],1007'd0},p_prime[1007],c_w_1007);
AND_array_1509 AND_array_1509_s1007({a_s[501:0],1007'd0},p_prime[1007],s_w_1007);
AND_array_1509 AND_array_1509_c1008({a_c[500:0],1008'd0},p_prime[1008],c_w_1008);
AND_array_1509 AND_array_1509_s1008({a_s[500:0],1008'd0},p_prime[1008],s_w_1008);
AND_array_1509 AND_array_1509_c1009({a_c[499:0],1009'd0},p_prime[1009],c_w_1009);
AND_array_1509 AND_array_1509_s1009({a_s[499:0],1009'd0},p_prime[1009],s_w_1009);
AND_array_1509 AND_array_1509_c1010({a_c[498:0],1010'd0},p_prime[1010],c_w_1010);
AND_array_1509 AND_array_1509_s1010({a_s[498:0],1010'd0},p_prime[1010],s_w_1010);
AND_array_1509 AND_array_1509_c1011({a_c[497:0],1011'd0},p_prime[1011],c_w_1011);
AND_array_1509 AND_array_1509_s1011({a_s[497:0],1011'd0},p_prime[1011],s_w_1011);
AND_array_1509 AND_array_1509_c1012({a_c[496:0],1012'd0},p_prime[1012],c_w_1012);
AND_array_1509 AND_array_1509_s1012({a_s[496:0],1012'd0},p_prime[1012],s_w_1012);
AND_array_1509 AND_array_1509_c1013({a_c[495:0],1013'd0},p_prime[1013],c_w_1013);
AND_array_1509 AND_array_1509_s1013({a_s[495:0],1013'd0},p_prime[1013],s_w_1013);
AND_array_1509 AND_array_1509_c1014({a_c[494:0],1014'd0},p_prime[1014],c_w_1014);
AND_array_1509 AND_array_1509_s1014({a_s[494:0],1014'd0},p_prime[1014],s_w_1014);
AND_array_1509 AND_array_1509_c1015({a_c[493:0],1015'd0},p_prime[1015],c_w_1015);
AND_array_1509 AND_array_1509_s1015({a_s[493:0],1015'd0},p_prime[1015],s_w_1015);
AND_array_1509 AND_array_1509_c1016({a_c[492:0],1016'd0},p_prime[1016],c_w_1016);
AND_array_1509 AND_array_1509_s1016({a_s[492:0],1016'd0},p_prime[1016],s_w_1016);
AND_array_1509 AND_array_1509_c1017({a_c[491:0],1017'd0},p_prime[1017],c_w_1017);
AND_array_1509 AND_array_1509_s1017({a_s[491:0],1017'd0},p_prime[1017],s_w_1017);
AND_array_1509 AND_array_1509_c1018({a_c[490:0],1018'd0},p_prime[1018],c_w_1018);
AND_array_1509 AND_array_1509_s1018({a_s[490:0],1018'd0},p_prime[1018],s_w_1018);
AND_array_1509 AND_array_1509_c1019({a_c[489:0],1019'd0},p_prime[1019],c_w_1019);
AND_array_1509 AND_array_1509_s1019({a_s[489:0],1019'd0},p_prime[1019],s_w_1019);
AND_array_1509 AND_array_1509_c1020({a_c[488:0],1020'd0},p_prime[1020],c_w_1020);
AND_array_1509 AND_array_1509_s1020({a_s[488:0],1020'd0},p_prime[1020],s_w_1020);
AND_array_1509 AND_array_1509_c1021({a_c[487:0],1021'd0},p_prime[1021],c_w_1021);
AND_array_1509 AND_array_1509_s1021({a_s[487:0],1021'd0},p_prime[1021],s_w_1021);
AND_array_1509 AND_array_1509_c1022({a_c[486:0],1022'd0},p_prime[1022],c_w_1022);
AND_array_1509 AND_array_1509_s1022({a_s[486:0],1022'd0},p_prime[1022],s_w_1022);
AND_array_1509 AND_array_1509_c1023({a_c[485:0],1023'd0},p_prime[1023],c_w_1023);
AND_array_1509 AND_array_1509_s1023({a_s[485:0],1023'd0},p_prime[1023],s_w_1023);
AND_array_1509 AND_array_1509_c1024({a_c[484:0],1024'd0},p_prime[1024],c_w_1024);
AND_array_1509 AND_array_1509_s1024({a_s[484:0],1024'd0},p_prime[1024],s_w_1024);
AND_array_1509 AND_array_1509_c1025({a_c[483:0],1025'd0},p_prime[1025],c_w_1025);
AND_array_1509 AND_array_1509_s1025({a_s[483:0],1025'd0},p_prime[1025],s_w_1025);
AND_array_1509 AND_array_1509_c1026({a_c[482:0],1026'd0},p_prime[1026],c_w_1026);
AND_array_1509 AND_array_1509_s1026({a_s[482:0],1026'd0},p_prime[1026],s_w_1026);
AND_array_1509 AND_array_1509_c1027({a_c[481:0],1027'd0},p_prime[1027],c_w_1027);
AND_array_1509 AND_array_1509_s1027({a_s[481:0],1027'd0},p_prime[1027],s_w_1027);
AND_array_1509 AND_array_1509_c1028({a_c[480:0],1028'd0},p_prime[1028],c_w_1028);
AND_array_1509 AND_array_1509_s1028({a_s[480:0],1028'd0},p_prime[1028],s_w_1028);
AND_array_1509 AND_array_1509_c1029({a_c[479:0],1029'd0},p_prime[1029],c_w_1029);
AND_array_1509 AND_array_1509_s1029({a_s[479:0],1029'd0},p_prime[1029],s_w_1029);
AND_array_1509 AND_array_1509_c1030({a_c[478:0],1030'd0},p_prime[1030],c_w_1030);
AND_array_1509 AND_array_1509_s1030({a_s[478:0],1030'd0},p_prime[1030],s_w_1030);
AND_array_1509 AND_array_1509_c1031({a_c[477:0],1031'd0},p_prime[1031],c_w_1031);
AND_array_1509 AND_array_1509_s1031({a_s[477:0],1031'd0},p_prime[1031],s_w_1031);
AND_array_1509 AND_array_1509_c1032({a_c[476:0],1032'd0},p_prime[1032],c_w_1032);
AND_array_1509 AND_array_1509_s1032({a_s[476:0],1032'd0},p_prime[1032],s_w_1032);
AND_array_1509 AND_array_1509_c1033({a_c[475:0],1033'd0},p_prime[1033],c_w_1033);
AND_array_1509 AND_array_1509_s1033({a_s[475:0],1033'd0},p_prime[1033],s_w_1033);
AND_array_1509 AND_array_1509_c1034({a_c[474:0],1034'd0},p_prime[1034],c_w_1034);
AND_array_1509 AND_array_1509_s1034({a_s[474:0],1034'd0},p_prime[1034],s_w_1034);
AND_array_1509 AND_array_1509_c1035({a_c[473:0],1035'd0},p_prime[1035],c_w_1035);
AND_array_1509 AND_array_1509_s1035({a_s[473:0],1035'd0},p_prime[1035],s_w_1035);
AND_array_1509 AND_array_1509_c1036({a_c[472:0],1036'd0},p_prime[1036],c_w_1036);
AND_array_1509 AND_array_1509_s1036({a_s[472:0],1036'd0},p_prime[1036],s_w_1036);
AND_array_1509 AND_array_1509_c1037({a_c[471:0],1037'd0},p_prime[1037],c_w_1037);
AND_array_1509 AND_array_1509_s1037({a_s[471:0],1037'd0},p_prime[1037],s_w_1037);
AND_array_1509 AND_array_1509_c1038({a_c[470:0],1038'd0},p_prime[1038],c_w_1038);
AND_array_1509 AND_array_1509_s1038({a_s[470:0],1038'd0},p_prime[1038],s_w_1038);
AND_array_1509 AND_array_1509_c1039({a_c[469:0],1039'd0},p_prime[1039],c_w_1039);
AND_array_1509 AND_array_1509_s1039({a_s[469:0],1039'd0},p_prime[1039],s_w_1039);
AND_array_1509 AND_array_1509_c1040({a_c[468:0],1040'd0},p_prime[1040],c_w_1040);
AND_array_1509 AND_array_1509_s1040({a_s[468:0],1040'd0},p_prime[1040],s_w_1040);
AND_array_1509 AND_array_1509_c1041({a_c[467:0],1041'd0},p_prime[1041],c_w_1041);
AND_array_1509 AND_array_1509_s1041({a_s[467:0],1041'd0},p_prime[1041],s_w_1041);
AND_array_1509 AND_array_1509_c1042({a_c[466:0],1042'd0},p_prime[1042],c_w_1042);
AND_array_1509 AND_array_1509_s1042({a_s[466:0],1042'd0},p_prime[1042],s_w_1042);
AND_array_1509 AND_array_1509_c1043({a_c[465:0],1043'd0},p_prime[1043],c_w_1043);
AND_array_1509 AND_array_1509_s1043({a_s[465:0],1043'd0},p_prime[1043],s_w_1043);
AND_array_1509 AND_array_1509_c1044({a_c[464:0],1044'd0},p_prime[1044],c_w_1044);
AND_array_1509 AND_array_1509_s1044({a_s[464:0],1044'd0},p_prime[1044],s_w_1044);
AND_array_1509 AND_array_1509_c1045({a_c[463:0],1045'd0},p_prime[1045],c_w_1045);
AND_array_1509 AND_array_1509_s1045({a_s[463:0],1045'd0},p_prime[1045],s_w_1045);
AND_array_1509 AND_array_1509_c1046({a_c[462:0],1046'd0},p_prime[1046],c_w_1046);
AND_array_1509 AND_array_1509_s1046({a_s[462:0],1046'd0},p_prime[1046],s_w_1046);
AND_array_1509 AND_array_1509_c1047({a_c[461:0],1047'd0},p_prime[1047],c_w_1047);
AND_array_1509 AND_array_1509_s1047({a_s[461:0],1047'd0},p_prime[1047],s_w_1047);
AND_array_1509 AND_array_1509_c1048({a_c[460:0],1048'd0},p_prime[1048],c_w_1048);
AND_array_1509 AND_array_1509_s1048({a_s[460:0],1048'd0},p_prime[1048],s_w_1048);
AND_array_1509 AND_array_1509_c1049({a_c[459:0],1049'd0},p_prime[1049],c_w_1049);
AND_array_1509 AND_array_1509_s1049({a_s[459:0],1049'd0},p_prime[1049],s_w_1049);
AND_array_1509 AND_array_1509_c1050({a_c[458:0],1050'd0},p_prime[1050],c_w_1050);
AND_array_1509 AND_array_1509_s1050({a_s[458:0],1050'd0},p_prime[1050],s_w_1050);
AND_array_1509 AND_array_1509_c1051({a_c[457:0],1051'd0},p_prime[1051],c_w_1051);
AND_array_1509 AND_array_1509_s1051({a_s[457:0],1051'd0},p_prime[1051],s_w_1051);
AND_array_1509 AND_array_1509_c1052({a_c[456:0],1052'd0},p_prime[1052],c_w_1052);
AND_array_1509 AND_array_1509_s1052({a_s[456:0],1052'd0},p_prime[1052],s_w_1052);
AND_array_1509 AND_array_1509_c1053({a_c[455:0],1053'd0},p_prime[1053],c_w_1053);
AND_array_1509 AND_array_1509_s1053({a_s[455:0],1053'd0},p_prime[1053],s_w_1053);
AND_array_1509 AND_array_1509_c1054({a_c[454:0],1054'd0},p_prime[1054],c_w_1054);
AND_array_1509 AND_array_1509_s1054({a_s[454:0],1054'd0},p_prime[1054],s_w_1054);
AND_array_1509 AND_array_1509_c1055({a_c[453:0],1055'd0},p_prime[1055],c_w_1055);
AND_array_1509 AND_array_1509_s1055({a_s[453:0],1055'd0},p_prime[1055],s_w_1055);
AND_array_1509 AND_array_1509_c1056({a_c[452:0],1056'd0},p_prime[1056],c_w_1056);
AND_array_1509 AND_array_1509_s1056({a_s[452:0],1056'd0},p_prime[1056],s_w_1056);
AND_array_1509 AND_array_1509_c1057({a_c[451:0],1057'd0},p_prime[1057],c_w_1057);
AND_array_1509 AND_array_1509_s1057({a_s[451:0],1057'd0},p_prime[1057],s_w_1057);
AND_array_1509 AND_array_1509_c1058({a_c[450:0],1058'd0},p_prime[1058],c_w_1058);
AND_array_1509 AND_array_1509_s1058({a_s[450:0],1058'd0},p_prime[1058],s_w_1058);
AND_array_1509 AND_array_1509_c1059({a_c[449:0],1059'd0},p_prime[1059],c_w_1059);
AND_array_1509 AND_array_1509_s1059({a_s[449:0],1059'd0},p_prime[1059],s_w_1059);
AND_array_1509 AND_array_1509_c1060({a_c[448:0],1060'd0},p_prime[1060],c_w_1060);
AND_array_1509 AND_array_1509_s1060({a_s[448:0],1060'd0},p_prime[1060],s_w_1060);
AND_array_1509 AND_array_1509_c1061({a_c[447:0],1061'd0},p_prime[1061],c_w_1061);
AND_array_1509 AND_array_1509_s1061({a_s[447:0],1061'd0},p_prime[1061],s_w_1061);
AND_array_1509 AND_array_1509_c1062({a_c[446:0],1062'd0},p_prime[1062],c_w_1062);
AND_array_1509 AND_array_1509_s1062({a_s[446:0],1062'd0},p_prime[1062],s_w_1062);
AND_array_1509 AND_array_1509_c1063({a_c[445:0],1063'd0},p_prime[1063],c_w_1063);
AND_array_1509 AND_array_1509_s1063({a_s[445:0],1063'd0},p_prime[1063],s_w_1063);
AND_array_1509 AND_array_1509_c1064({a_c[444:0],1064'd0},p_prime[1064],c_w_1064);
AND_array_1509 AND_array_1509_s1064({a_s[444:0],1064'd0},p_prime[1064],s_w_1064);
AND_array_1509 AND_array_1509_c1065({a_c[443:0],1065'd0},p_prime[1065],c_w_1065);
AND_array_1509 AND_array_1509_s1065({a_s[443:0],1065'd0},p_prime[1065],s_w_1065);
AND_array_1509 AND_array_1509_c1066({a_c[442:0],1066'd0},p_prime[1066],c_w_1066);
AND_array_1509 AND_array_1509_s1066({a_s[442:0],1066'd0},p_prime[1066],s_w_1066);
AND_array_1509 AND_array_1509_c1067({a_c[441:0],1067'd0},p_prime[1067],c_w_1067);
AND_array_1509 AND_array_1509_s1067({a_s[441:0],1067'd0},p_prime[1067],s_w_1067);
AND_array_1509 AND_array_1509_c1068({a_c[440:0],1068'd0},p_prime[1068],c_w_1068);
AND_array_1509 AND_array_1509_s1068({a_s[440:0],1068'd0},p_prime[1068],s_w_1068);
AND_array_1509 AND_array_1509_c1069({a_c[439:0],1069'd0},p_prime[1069],c_w_1069);
AND_array_1509 AND_array_1509_s1069({a_s[439:0],1069'd0},p_prime[1069],s_w_1069);
AND_array_1509 AND_array_1509_c1070({a_c[438:0],1070'd0},p_prime[1070],c_w_1070);
AND_array_1509 AND_array_1509_s1070({a_s[438:0],1070'd0},p_prime[1070],s_w_1070);
AND_array_1509 AND_array_1509_c1071({a_c[437:0],1071'd0},p_prime[1071],c_w_1071);
AND_array_1509 AND_array_1509_s1071({a_s[437:0],1071'd0},p_prime[1071],s_w_1071);
AND_array_1509 AND_array_1509_c1072({a_c[436:0],1072'd0},p_prime[1072],c_w_1072);
AND_array_1509 AND_array_1509_s1072({a_s[436:0],1072'd0},p_prime[1072],s_w_1072);
AND_array_1509 AND_array_1509_c1073({a_c[435:0],1073'd0},p_prime[1073],c_w_1073);
AND_array_1509 AND_array_1509_s1073({a_s[435:0],1073'd0},p_prime[1073],s_w_1073);
AND_array_1509 AND_array_1509_c1074({a_c[434:0],1074'd0},p_prime[1074],c_w_1074);
AND_array_1509 AND_array_1509_s1074({a_s[434:0],1074'd0},p_prime[1074],s_w_1074);
AND_array_1509 AND_array_1509_c1075({a_c[433:0],1075'd0},p_prime[1075],c_w_1075);
AND_array_1509 AND_array_1509_s1075({a_s[433:0],1075'd0},p_prime[1075],s_w_1075);
AND_array_1509 AND_array_1509_c1076({a_c[432:0],1076'd0},p_prime[1076],c_w_1076);
AND_array_1509 AND_array_1509_s1076({a_s[432:0],1076'd0},p_prime[1076],s_w_1076);
AND_array_1509 AND_array_1509_c1077({a_c[431:0],1077'd0},p_prime[1077],c_w_1077);
AND_array_1509 AND_array_1509_s1077({a_s[431:0],1077'd0},p_prime[1077],s_w_1077);
AND_array_1509 AND_array_1509_c1078({a_c[430:0],1078'd0},p_prime[1078],c_w_1078);
AND_array_1509 AND_array_1509_s1078({a_s[430:0],1078'd0},p_prime[1078],s_w_1078);
AND_array_1509 AND_array_1509_c1079({a_c[429:0],1079'd0},p_prime[1079],c_w_1079);
AND_array_1509 AND_array_1509_s1079({a_s[429:0],1079'd0},p_prime[1079],s_w_1079);
AND_array_1509 AND_array_1509_c1080({a_c[428:0],1080'd0},p_prime[1080],c_w_1080);
AND_array_1509 AND_array_1509_s1080({a_s[428:0],1080'd0},p_prime[1080],s_w_1080);
AND_array_1509 AND_array_1509_c1081({a_c[427:0],1081'd0},p_prime[1081],c_w_1081);
AND_array_1509 AND_array_1509_s1081({a_s[427:0],1081'd0},p_prime[1081],s_w_1081);
AND_array_1509 AND_array_1509_c1082({a_c[426:0],1082'd0},p_prime[1082],c_w_1082);
AND_array_1509 AND_array_1509_s1082({a_s[426:0],1082'd0},p_prime[1082],s_w_1082);
AND_array_1509 AND_array_1509_c1083({a_c[425:0],1083'd0},p_prime[1083],c_w_1083);
AND_array_1509 AND_array_1509_s1083({a_s[425:0],1083'd0},p_prime[1083],s_w_1083);
AND_array_1509 AND_array_1509_c1084({a_c[424:0],1084'd0},p_prime[1084],c_w_1084);
AND_array_1509 AND_array_1509_s1084({a_s[424:0],1084'd0},p_prime[1084],s_w_1084);
AND_array_1509 AND_array_1509_c1085({a_c[423:0],1085'd0},p_prime[1085],c_w_1085);
AND_array_1509 AND_array_1509_s1085({a_s[423:0],1085'd0},p_prime[1085],s_w_1085);
AND_array_1509 AND_array_1509_c1086({a_c[422:0],1086'd0},p_prime[1086],c_w_1086);
AND_array_1509 AND_array_1509_s1086({a_s[422:0],1086'd0},p_prime[1086],s_w_1086);
AND_array_1509 AND_array_1509_c1087({a_c[421:0],1087'd0},p_prime[1087],c_w_1087);
AND_array_1509 AND_array_1509_s1087({a_s[421:0],1087'd0},p_prime[1087],s_w_1087);
AND_array_1509 AND_array_1509_c1088({a_c[420:0],1088'd0},p_prime[1088],c_w_1088);
AND_array_1509 AND_array_1509_s1088({a_s[420:0],1088'd0},p_prime[1088],s_w_1088);
AND_array_1509 AND_array_1509_c1089({a_c[419:0],1089'd0},p_prime[1089],c_w_1089);
AND_array_1509 AND_array_1509_s1089({a_s[419:0],1089'd0},p_prime[1089],s_w_1089);
AND_array_1509 AND_array_1509_c1090({a_c[418:0],1090'd0},p_prime[1090],c_w_1090);
AND_array_1509 AND_array_1509_s1090({a_s[418:0],1090'd0},p_prime[1090],s_w_1090);
AND_array_1509 AND_array_1509_c1091({a_c[417:0],1091'd0},p_prime[1091],c_w_1091);
AND_array_1509 AND_array_1509_s1091({a_s[417:0],1091'd0},p_prime[1091],s_w_1091);
AND_array_1509 AND_array_1509_c1092({a_c[416:0],1092'd0},p_prime[1092],c_w_1092);
AND_array_1509 AND_array_1509_s1092({a_s[416:0],1092'd0},p_prime[1092],s_w_1092);
AND_array_1509 AND_array_1509_c1093({a_c[415:0],1093'd0},p_prime[1093],c_w_1093);
AND_array_1509 AND_array_1509_s1093({a_s[415:0],1093'd0},p_prime[1093],s_w_1093);
AND_array_1509 AND_array_1509_c1094({a_c[414:0],1094'd0},p_prime[1094],c_w_1094);
AND_array_1509 AND_array_1509_s1094({a_s[414:0],1094'd0},p_prime[1094],s_w_1094);
AND_array_1509 AND_array_1509_c1095({a_c[413:0],1095'd0},p_prime[1095],c_w_1095);
AND_array_1509 AND_array_1509_s1095({a_s[413:0],1095'd0},p_prime[1095],s_w_1095);
AND_array_1509 AND_array_1509_c1096({a_c[412:0],1096'd0},p_prime[1096],c_w_1096);
AND_array_1509 AND_array_1509_s1096({a_s[412:0],1096'd0},p_prime[1096],s_w_1096);
AND_array_1509 AND_array_1509_c1097({a_c[411:0],1097'd0},p_prime[1097],c_w_1097);
AND_array_1509 AND_array_1509_s1097({a_s[411:0],1097'd0},p_prime[1097],s_w_1097);
AND_array_1509 AND_array_1509_c1098({a_c[410:0],1098'd0},p_prime[1098],c_w_1098);
AND_array_1509 AND_array_1509_s1098({a_s[410:0],1098'd0},p_prime[1098],s_w_1098);
AND_array_1509 AND_array_1509_c1099({a_c[409:0],1099'd0},p_prime[1099],c_w_1099);
AND_array_1509 AND_array_1509_s1099({a_s[409:0],1099'd0},p_prime[1099],s_w_1099);
AND_array_1509 AND_array_1509_c1100({a_c[408:0],1100'd0},p_prime[1100],c_w_1100);
AND_array_1509 AND_array_1509_s1100({a_s[408:0],1100'd0},p_prime[1100],s_w_1100);
AND_array_1509 AND_array_1509_c1101({a_c[407:0],1101'd0},p_prime[1101],c_w_1101);
AND_array_1509 AND_array_1509_s1101({a_s[407:0],1101'd0},p_prime[1101],s_w_1101);
AND_array_1509 AND_array_1509_c1102({a_c[406:0],1102'd0},p_prime[1102],c_w_1102);
AND_array_1509 AND_array_1509_s1102({a_s[406:0],1102'd0},p_prime[1102],s_w_1102);
AND_array_1509 AND_array_1509_c1103({a_c[405:0],1103'd0},p_prime[1103],c_w_1103);
AND_array_1509 AND_array_1509_s1103({a_s[405:0],1103'd0},p_prime[1103],s_w_1103);
AND_array_1509 AND_array_1509_c1104({a_c[404:0],1104'd0},p_prime[1104],c_w_1104);
AND_array_1509 AND_array_1509_s1104({a_s[404:0],1104'd0},p_prime[1104],s_w_1104);
AND_array_1509 AND_array_1509_c1105({a_c[403:0],1105'd0},p_prime[1105],c_w_1105);
AND_array_1509 AND_array_1509_s1105({a_s[403:0],1105'd0},p_prime[1105],s_w_1105);
AND_array_1509 AND_array_1509_c1106({a_c[402:0],1106'd0},p_prime[1106],c_w_1106);
AND_array_1509 AND_array_1509_s1106({a_s[402:0],1106'd0},p_prime[1106],s_w_1106);
AND_array_1509 AND_array_1509_c1107({a_c[401:0],1107'd0},p_prime[1107],c_w_1107);
AND_array_1509 AND_array_1509_s1107({a_s[401:0],1107'd0},p_prime[1107],s_w_1107);
AND_array_1509 AND_array_1509_c1108({a_c[400:0],1108'd0},p_prime[1108],c_w_1108);
AND_array_1509 AND_array_1509_s1108({a_s[400:0],1108'd0},p_prime[1108],s_w_1108);
AND_array_1509 AND_array_1509_c1109({a_c[399:0],1109'd0},p_prime[1109],c_w_1109);
AND_array_1509 AND_array_1509_s1109({a_s[399:0],1109'd0},p_prime[1109],s_w_1109);
AND_array_1509 AND_array_1509_c1110({a_c[398:0],1110'd0},p_prime[1110],c_w_1110);
AND_array_1509 AND_array_1509_s1110({a_s[398:0],1110'd0},p_prime[1110],s_w_1110);
AND_array_1509 AND_array_1509_c1111({a_c[397:0],1111'd0},p_prime[1111],c_w_1111);
AND_array_1509 AND_array_1509_s1111({a_s[397:0],1111'd0},p_prime[1111],s_w_1111);
AND_array_1509 AND_array_1509_c1112({a_c[396:0],1112'd0},p_prime[1112],c_w_1112);
AND_array_1509 AND_array_1509_s1112({a_s[396:0],1112'd0},p_prime[1112],s_w_1112);
AND_array_1509 AND_array_1509_c1113({a_c[395:0],1113'd0},p_prime[1113],c_w_1113);
AND_array_1509 AND_array_1509_s1113({a_s[395:0],1113'd0},p_prime[1113],s_w_1113);
AND_array_1509 AND_array_1509_c1114({a_c[394:0],1114'd0},p_prime[1114],c_w_1114);
AND_array_1509 AND_array_1509_s1114({a_s[394:0],1114'd0},p_prime[1114],s_w_1114);
AND_array_1509 AND_array_1509_c1115({a_c[393:0],1115'd0},p_prime[1115],c_w_1115);
AND_array_1509 AND_array_1509_s1115({a_s[393:0],1115'd0},p_prime[1115],s_w_1115);
AND_array_1509 AND_array_1509_c1116({a_c[392:0],1116'd0},p_prime[1116],c_w_1116);
AND_array_1509 AND_array_1509_s1116({a_s[392:0],1116'd0},p_prime[1116],s_w_1116);
AND_array_1509 AND_array_1509_c1117({a_c[391:0],1117'd0},p_prime[1117],c_w_1117);
AND_array_1509 AND_array_1509_s1117({a_s[391:0],1117'd0},p_prime[1117],s_w_1117);
AND_array_1509 AND_array_1509_c1118({a_c[390:0],1118'd0},p_prime[1118],c_w_1118);
AND_array_1509 AND_array_1509_s1118({a_s[390:0],1118'd0},p_prime[1118],s_w_1118);
AND_array_1509 AND_array_1509_c1119({a_c[389:0],1119'd0},p_prime[1119],c_w_1119);
AND_array_1509 AND_array_1509_s1119({a_s[389:0],1119'd0},p_prime[1119],s_w_1119);
AND_array_1509 AND_array_1509_c1120({a_c[388:0],1120'd0},p_prime[1120],c_w_1120);
AND_array_1509 AND_array_1509_s1120({a_s[388:0],1120'd0},p_prime[1120],s_w_1120);
AND_array_1509 AND_array_1509_c1121({a_c[387:0],1121'd0},p_prime[1121],c_w_1121);
AND_array_1509 AND_array_1509_s1121({a_s[387:0],1121'd0},p_prime[1121],s_w_1121);
AND_array_1509 AND_array_1509_c1122({a_c[386:0],1122'd0},p_prime[1122],c_w_1122);
AND_array_1509 AND_array_1509_s1122({a_s[386:0],1122'd0},p_prime[1122],s_w_1122);
AND_array_1509 AND_array_1509_c1123({a_c[385:0],1123'd0},p_prime[1123],c_w_1123);
AND_array_1509 AND_array_1509_s1123({a_s[385:0],1123'd0},p_prime[1123],s_w_1123);
AND_array_1509 AND_array_1509_c1124({a_c[384:0],1124'd0},p_prime[1124],c_w_1124);
AND_array_1509 AND_array_1509_s1124({a_s[384:0],1124'd0},p_prime[1124],s_w_1124);
AND_array_1509 AND_array_1509_c1125({a_c[383:0],1125'd0},p_prime[1125],c_w_1125);
AND_array_1509 AND_array_1509_s1125({a_s[383:0],1125'd0},p_prime[1125],s_w_1125);
AND_array_1509 AND_array_1509_c1126({a_c[382:0],1126'd0},p_prime[1126],c_w_1126);
AND_array_1509 AND_array_1509_s1126({a_s[382:0],1126'd0},p_prime[1126],s_w_1126);
AND_array_1509 AND_array_1509_c1127({a_c[381:0],1127'd0},p_prime[1127],c_w_1127);
AND_array_1509 AND_array_1509_s1127({a_s[381:0],1127'd0},p_prime[1127],s_w_1127);
AND_array_1509 AND_array_1509_c1128({a_c[380:0],1128'd0},p_prime[1128],c_w_1128);
AND_array_1509 AND_array_1509_s1128({a_s[380:0],1128'd0},p_prime[1128],s_w_1128);
AND_array_1509 AND_array_1509_c1129({a_c[379:0],1129'd0},p_prime[1129],c_w_1129);
AND_array_1509 AND_array_1509_s1129({a_s[379:0],1129'd0},p_prime[1129],s_w_1129);
AND_array_1509 AND_array_1509_c1130({a_c[378:0],1130'd0},p_prime[1130],c_w_1130);
AND_array_1509 AND_array_1509_s1130({a_s[378:0],1130'd0},p_prime[1130],s_w_1130);
AND_array_1509 AND_array_1509_c1131({a_c[377:0],1131'd0},p_prime[1131],c_w_1131);
AND_array_1509 AND_array_1509_s1131({a_s[377:0],1131'd0},p_prime[1131],s_w_1131);
AND_array_1509 AND_array_1509_c1132({a_c[376:0],1132'd0},p_prime[1132],c_w_1132);
AND_array_1509 AND_array_1509_s1132({a_s[376:0],1132'd0},p_prime[1132],s_w_1132);
AND_array_1509 AND_array_1509_c1133({a_c[375:0],1133'd0},p_prime[1133],c_w_1133);
AND_array_1509 AND_array_1509_s1133({a_s[375:0],1133'd0},p_prime[1133],s_w_1133);
AND_array_1509 AND_array_1509_c1134({a_c[374:0],1134'd0},p_prime[1134],c_w_1134);
AND_array_1509 AND_array_1509_s1134({a_s[374:0],1134'd0},p_prime[1134],s_w_1134);
AND_array_1509 AND_array_1509_c1135({a_c[373:0],1135'd0},p_prime[1135],c_w_1135);
AND_array_1509 AND_array_1509_s1135({a_s[373:0],1135'd0},p_prime[1135],s_w_1135);
AND_array_1509 AND_array_1509_c1136({a_c[372:0],1136'd0},p_prime[1136],c_w_1136);
AND_array_1509 AND_array_1509_s1136({a_s[372:0],1136'd0},p_prime[1136],s_w_1136);
AND_array_1509 AND_array_1509_c1137({a_c[371:0],1137'd0},p_prime[1137],c_w_1137);
AND_array_1509 AND_array_1509_s1137({a_s[371:0],1137'd0},p_prime[1137],s_w_1137);
AND_array_1509 AND_array_1509_c1138({a_c[370:0],1138'd0},p_prime[1138],c_w_1138);
AND_array_1509 AND_array_1509_s1138({a_s[370:0],1138'd0},p_prime[1138],s_w_1138);
AND_array_1509 AND_array_1509_c1139({a_c[369:0],1139'd0},p_prime[1139],c_w_1139);
AND_array_1509 AND_array_1509_s1139({a_s[369:0],1139'd0},p_prime[1139],s_w_1139);
AND_array_1509 AND_array_1509_c1140({a_c[368:0],1140'd0},p_prime[1140],c_w_1140);
AND_array_1509 AND_array_1509_s1140({a_s[368:0],1140'd0},p_prime[1140],s_w_1140);
AND_array_1509 AND_array_1509_c1141({a_c[367:0],1141'd0},p_prime[1141],c_w_1141);
AND_array_1509 AND_array_1509_s1141({a_s[367:0],1141'd0},p_prime[1141],s_w_1141);
AND_array_1509 AND_array_1509_c1142({a_c[366:0],1142'd0},p_prime[1142],c_w_1142);
AND_array_1509 AND_array_1509_s1142({a_s[366:0],1142'd0},p_prime[1142],s_w_1142);
AND_array_1509 AND_array_1509_c1143({a_c[365:0],1143'd0},p_prime[1143],c_w_1143);
AND_array_1509 AND_array_1509_s1143({a_s[365:0],1143'd0},p_prime[1143],s_w_1143);
AND_array_1509 AND_array_1509_c1144({a_c[364:0],1144'd0},p_prime[1144],c_w_1144);
AND_array_1509 AND_array_1509_s1144({a_s[364:0],1144'd0},p_prime[1144],s_w_1144);
AND_array_1509 AND_array_1509_c1145({a_c[363:0],1145'd0},p_prime[1145],c_w_1145);
AND_array_1509 AND_array_1509_s1145({a_s[363:0],1145'd0},p_prime[1145],s_w_1145);
AND_array_1509 AND_array_1509_c1146({a_c[362:0],1146'd0},p_prime[1146],c_w_1146);
AND_array_1509 AND_array_1509_s1146({a_s[362:0],1146'd0},p_prime[1146],s_w_1146);
AND_array_1509 AND_array_1509_c1147({a_c[361:0],1147'd0},p_prime[1147],c_w_1147);
AND_array_1509 AND_array_1509_s1147({a_s[361:0],1147'd0},p_prime[1147],s_w_1147);
AND_array_1509 AND_array_1509_c1148({a_c[360:0],1148'd0},p_prime[1148],c_w_1148);
AND_array_1509 AND_array_1509_s1148({a_s[360:0],1148'd0},p_prime[1148],s_w_1148);
AND_array_1509 AND_array_1509_c1149({a_c[359:0],1149'd0},p_prime[1149],c_w_1149);
AND_array_1509 AND_array_1509_s1149({a_s[359:0],1149'd0},p_prime[1149],s_w_1149);
AND_array_1509 AND_array_1509_c1150({a_c[358:0],1150'd0},p_prime[1150],c_w_1150);
AND_array_1509 AND_array_1509_s1150({a_s[358:0],1150'd0},p_prime[1150],s_w_1150);
AND_array_1509 AND_array_1509_c1151({a_c[357:0],1151'd0},p_prime[1151],c_w_1151);
AND_array_1509 AND_array_1509_s1151({a_s[357:0],1151'd0},p_prime[1151],s_w_1151);
AND_array_1509 AND_array_1509_c1152({a_c[356:0],1152'd0},p_prime[1152],c_w_1152);
AND_array_1509 AND_array_1509_s1152({a_s[356:0],1152'd0},p_prime[1152],s_w_1152);
AND_array_1509 AND_array_1509_c1153({a_c[355:0],1153'd0},p_prime[1153],c_w_1153);
AND_array_1509 AND_array_1509_s1153({a_s[355:0],1153'd0},p_prime[1153],s_w_1153);
AND_array_1509 AND_array_1509_c1154({a_c[354:0],1154'd0},p_prime[1154],c_w_1154);
AND_array_1509 AND_array_1509_s1154({a_s[354:0],1154'd0},p_prime[1154],s_w_1154);
AND_array_1509 AND_array_1509_c1155({a_c[353:0],1155'd0},p_prime[1155],c_w_1155);
AND_array_1509 AND_array_1509_s1155({a_s[353:0],1155'd0},p_prime[1155],s_w_1155);
AND_array_1509 AND_array_1509_c1156({a_c[352:0],1156'd0},p_prime[1156],c_w_1156);
AND_array_1509 AND_array_1509_s1156({a_s[352:0],1156'd0},p_prime[1156],s_w_1156);
AND_array_1509 AND_array_1509_c1157({a_c[351:0],1157'd0},p_prime[1157],c_w_1157);
AND_array_1509 AND_array_1509_s1157({a_s[351:0],1157'd0},p_prime[1157],s_w_1157);
AND_array_1509 AND_array_1509_c1158({a_c[350:0],1158'd0},p_prime[1158],c_w_1158);
AND_array_1509 AND_array_1509_s1158({a_s[350:0],1158'd0},p_prime[1158],s_w_1158);
AND_array_1509 AND_array_1509_c1159({a_c[349:0],1159'd0},p_prime[1159],c_w_1159);
AND_array_1509 AND_array_1509_s1159({a_s[349:0],1159'd0},p_prime[1159],s_w_1159);
AND_array_1509 AND_array_1509_c1160({a_c[348:0],1160'd0},p_prime[1160],c_w_1160);
AND_array_1509 AND_array_1509_s1160({a_s[348:0],1160'd0},p_prime[1160],s_w_1160);
AND_array_1509 AND_array_1509_c1161({a_c[347:0],1161'd0},p_prime[1161],c_w_1161);
AND_array_1509 AND_array_1509_s1161({a_s[347:0],1161'd0},p_prime[1161],s_w_1161);
AND_array_1509 AND_array_1509_c1162({a_c[346:0],1162'd0},p_prime[1162],c_w_1162);
AND_array_1509 AND_array_1509_s1162({a_s[346:0],1162'd0},p_prime[1162],s_w_1162);
AND_array_1509 AND_array_1509_c1163({a_c[345:0],1163'd0},p_prime[1163],c_w_1163);
AND_array_1509 AND_array_1509_s1163({a_s[345:0],1163'd0},p_prime[1163],s_w_1163);
AND_array_1509 AND_array_1509_c1164({a_c[344:0],1164'd0},p_prime[1164],c_w_1164);
AND_array_1509 AND_array_1509_s1164({a_s[344:0],1164'd0},p_prime[1164],s_w_1164);
AND_array_1509 AND_array_1509_c1165({a_c[343:0],1165'd0},p_prime[1165],c_w_1165);
AND_array_1509 AND_array_1509_s1165({a_s[343:0],1165'd0},p_prime[1165],s_w_1165);
AND_array_1509 AND_array_1509_c1166({a_c[342:0],1166'd0},p_prime[1166],c_w_1166);
AND_array_1509 AND_array_1509_s1166({a_s[342:0],1166'd0},p_prime[1166],s_w_1166);
AND_array_1509 AND_array_1509_c1167({a_c[341:0],1167'd0},p_prime[1167],c_w_1167);
AND_array_1509 AND_array_1509_s1167({a_s[341:0],1167'd0},p_prime[1167],s_w_1167);
AND_array_1509 AND_array_1509_c1168({a_c[340:0],1168'd0},p_prime[1168],c_w_1168);
AND_array_1509 AND_array_1509_s1168({a_s[340:0],1168'd0},p_prime[1168],s_w_1168);
AND_array_1509 AND_array_1509_c1169({a_c[339:0],1169'd0},p_prime[1169],c_w_1169);
AND_array_1509 AND_array_1509_s1169({a_s[339:0],1169'd0},p_prime[1169],s_w_1169);
AND_array_1509 AND_array_1509_c1170({a_c[338:0],1170'd0},p_prime[1170],c_w_1170);
AND_array_1509 AND_array_1509_s1170({a_s[338:0],1170'd0},p_prime[1170],s_w_1170);
AND_array_1509 AND_array_1509_c1171({a_c[337:0],1171'd0},p_prime[1171],c_w_1171);
AND_array_1509 AND_array_1509_s1171({a_s[337:0],1171'd0},p_prime[1171],s_w_1171);
AND_array_1509 AND_array_1509_c1172({a_c[336:0],1172'd0},p_prime[1172],c_w_1172);
AND_array_1509 AND_array_1509_s1172({a_s[336:0],1172'd0},p_prime[1172],s_w_1172);
AND_array_1509 AND_array_1509_c1173({a_c[335:0],1173'd0},p_prime[1173],c_w_1173);
AND_array_1509 AND_array_1509_s1173({a_s[335:0],1173'd0},p_prime[1173],s_w_1173);
AND_array_1509 AND_array_1509_c1174({a_c[334:0],1174'd0},p_prime[1174],c_w_1174);
AND_array_1509 AND_array_1509_s1174({a_s[334:0],1174'd0},p_prime[1174],s_w_1174);
AND_array_1509 AND_array_1509_c1175({a_c[333:0],1175'd0},p_prime[1175],c_w_1175);
AND_array_1509 AND_array_1509_s1175({a_s[333:0],1175'd0},p_prime[1175],s_w_1175);
AND_array_1509 AND_array_1509_c1176({a_c[332:0],1176'd0},p_prime[1176],c_w_1176);
AND_array_1509 AND_array_1509_s1176({a_s[332:0],1176'd0},p_prime[1176],s_w_1176);
AND_array_1509 AND_array_1509_c1177({a_c[331:0],1177'd0},p_prime[1177],c_w_1177);
AND_array_1509 AND_array_1509_s1177({a_s[331:0],1177'd0},p_prime[1177],s_w_1177);
AND_array_1509 AND_array_1509_c1178({a_c[330:0],1178'd0},p_prime[1178],c_w_1178);
AND_array_1509 AND_array_1509_s1178({a_s[330:0],1178'd0},p_prime[1178],s_w_1178);
AND_array_1509 AND_array_1509_c1179({a_c[329:0],1179'd0},p_prime[1179],c_w_1179);
AND_array_1509 AND_array_1509_s1179({a_s[329:0],1179'd0},p_prime[1179],s_w_1179);
AND_array_1509 AND_array_1509_c1180({a_c[328:0],1180'd0},p_prime[1180],c_w_1180);
AND_array_1509 AND_array_1509_s1180({a_s[328:0],1180'd0},p_prime[1180],s_w_1180);
AND_array_1509 AND_array_1509_c1181({a_c[327:0],1181'd0},p_prime[1181],c_w_1181);
AND_array_1509 AND_array_1509_s1181({a_s[327:0],1181'd0},p_prime[1181],s_w_1181);
AND_array_1509 AND_array_1509_c1182({a_c[326:0],1182'd0},p_prime[1182],c_w_1182);
AND_array_1509 AND_array_1509_s1182({a_s[326:0],1182'd0},p_prime[1182],s_w_1182);
AND_array_1509 AND_array_1509_c1183({a_c[325:0],1183'd0},p_prime[1183],c_w_1183);
AND_array_1509 AND_array_1509_s1183({a_s[325:0],1183'd0},p_prime[1183],s_w_1183);
AND_array_1509 AND_array_1509_c1184({a_c[324:0],1184'd0},p_prime[1184],c_w_1184);
AND_array_1509 AND_array_1509_s1184({a_s[324:0],1184'd0},p_prime[1184],s_w_1184);
AND_array_1509 AND_array_1509_c1185({a_c[323:0],1185'd0},p_prime[1185],c_w_1185);
AND_array_1509 AND_array_1509_s1185({a_s[323:0],1185'd0},p_prime[1185],s_w_1185);
AND_array_1509 AND_array_1509_c1186({a_c[322:0],1186'd0},p_prime[1186],c_w_1186);
AND_array_1509 AND_array_1509_s1186({a_s[322:0],1186'd0},p_prime[1186],s_w_1186);
AND_array_1509 AND_array_1509_c1187({a_c[321:0],1187'd0},p_prime[1187],c_w_1187);
AND_array_1509 AND_array_1509_s1187({a_s[321:0],1187'd0},p_prime[1187],s_w_1187);
AND_array_1509 AND_array_1509_c1188({a_c[320:0],1188'd0},p_prime[1188],c_w_1188);
AND_array_1509 AND_array_1509_s1188({a_s[320:0],1188'd0},p_prime[1188],s_w_1188);
AND_array_1509 AND_array_1509_c1189({a_c[319:0],1189'd0},p_prime[1189],c_w_1189);
AND_array_1509 AND_array_1509_s1189({a_s[319:0],1189'd0},p_prime[1189],s_w_1189);
AND_array_1509 AND_array_1509_c1190({a_c[318:0],1190'd0},p_prime[1190],c_w_1190);
AND_array_1509 AND_array_1509_s1190({a_s[318:0],1190'd0},p_prime[1190],s_w_1190);
AND_array_1509 AND_array_1509_c1191({a_c[317:0],1191'd0},p_prime[1191],c_w_1191);
AND_array_1509 AND_array_1509_s1191({a_s[317:0],1191'd0},p_prime[1191],s_w_1191);
AND_array_1509 AND_array_1509_c1192({a_c[316:0],1192'd0},p_prime[1192],c_w_1192);
AND_array_1509 AND_array_1509_s1192({a_s[316:0],1192'd0},p_prime[1192],s_w_1192);
AND_array_1509 AND_array_1509_c1193({a_c[315:0],1193'd0},p_prime[1193],c_w_1193);
AND_array_1509 AND_array_1509_s1193({a_s[315:0],1193'd0},p_prime[1193],s_w_1193);
AND_array_1509 AND_array_1509_c1194({a_c[314:0],1194'd0},p_prime[1194],c_w_1194);
AND_array_1509 AND_array_1509_s1194({a_s[314:0],1194'd0},p_prime[1194],s_w_1194);
AND_array_1509 AND_array_1509_c1195({a_c[313:0],1195'd0},p_prime[1195],c_w_1195);
AND_array_1509 AND_array_1509_s1195({a_s[313:0],1195'd0},p_prime[1195],s_w_1195);
AND_array_1509 AND_array_1509_c1196({a_c[312:0],1196'd0},p_prime[1196],c_w_1196);
AND_array_1509 AND_array_1509_s1196({a_s[312:0],1196'd0},p_prime[1196],s_w_1196);
AND_array_1509 AND_array_1509_c1197({a_c[311:0],1197'd0},p_prime[1197],c_w_1197);
AND_array_1509 AND_array_1509_s1197({a_s[311:0],1197'd0},p_prime[1197],s_w_1197);
AND_array_1509 AND_array_1509_c1198({a_c[310:0],1198'd0},p_prime[1198],c_w_1198);
AND_array_1509 AND_array_1509_s1198({a_s[310:0],1198'd0},p_prime[1198],s_w_1198);
AND_array_1509 AND_array_1509_c1199({a_c[309:0],1199'd0},p_prime[1199],c_w_1199);
AND_array_1509 AND_array_1509_s1199({a_s[309:0],1199'd0},p_prime[1199],s_w_1199);
AND_array_1509 AND_array_1509_c1200({a_c[308:0],1200'd0},p_prime[1200],c_w_1200);
AND_array_1509 AND_array_1509_s1200({a_s[308:0],1200'd0},p_prime[1200],s_w_1200);
AND_array_1509 AND_array_1509_c1201({a_c[307:0],1201'd0},p_prime[1201],c_w_1201);
AND_array_1509 AND_array_1509_s1201({a_s[307:0],1201'd0},p_prime[1201],s_w_1201);
AND_array_1509 AND_array_1509_c1202({a_c[306:0],1202'd0},p_prime[1202],c_w_1202);
AND_array_1509 AND_array_1509_s1202({a_s[306:0],1202'd0},p_prime[1202],s_w_1202);
AND_array_1509 AND_array_1509_c1203({a_c[305:0],1203'd0},p_prime[1203],c_w_1203);
AND_array_1509 AND_array_1509_s1203({a_s[305:0],1203'd0},p_prime[1203],s_w_1203);
AND_array_1509 AND_array_1509_c1204({a_c[304:0],1204'd0},p_prime[1204],c_w_1204);
AND_array_1509 AND_array_1509_s1204({a_s[304:0],1204'd0},p_prime[1204],s_w_1204);
AND_array_1509 AND_array_1509_c1205({a_c[303:0],1205'd0},p_prime[1205],c_w_1205);
AND_array_1509 AND_array_1509_s1205({a_s[303:0],1205'd0},p_prime[1205],s_w_1205);
AND_array_1509 AND_array_1509_c1206({a_c[302:0],1206'd0},p_prime[1206],c_w_1206);
AND_array_1509 AND_array_1509_s1206({a_s[302:0],1206'd0},p_prime[1206],s_w_1206);
AND_array_1509 AND_array_1509_c1207({a_c[301:0],1207'd0},p_prime[1207],c_w_1207);
AND_array_1509 AND_array_1509_s1207({a_s[301:0],1207'd0},p_prime[1207],s_w_1207);
AND_array_1509 AND_array_1509_c1208({a_c[300:0],1208'd0},p_prime[1208],c_w_1208);
AND_array_1509 AND_array_1509_s1208({a_s[300:0],1208'd0},p_prime[1208],s_w_1208);
AND_array_1509 AND_array_1509_c1209({a_c[299:0],1209'd0},p_prime[1209],c_w_1209);
AND_array_1509 AND_array_1509_s1209({a_s[299:0],1209'd0},p_prime[1209],s_w_1209);
AND_array_1509 AND_array_1509_c1210({a_c[298:0],1210'd0},p_prime[1210],c_w_1210);
AND_array_1509 AND_array_1509_s1210({a_s[298:0],1210'd0},p_prime[1210],s_w_1210);
AND_array_1509 AND_array_1509_c1211({a_c[297:0],1211'd0},p_prime[1211],c_w_1211);
AND_array_1509 AND_array_1509_s1211({a_s[297:0],1211'd0},p_prime[1211],s_w_1211);
AND_array_1509 AND_array_1509_c1212({a_c[296:0],1212'd0},p_prime[1212],c_w_1212);
AND_array_1509 AND_array_1509_s1212({a_s[296:0],1212'd0},p_prime[1212],s_w_1212);
AND_array_1509 AND_array_1509_c1213({a_c[295:0],1213'd0},p_prime[1213],c_w_1213);
AND_array_1509 AND_array_1509_s1213({a_s[295:0],1213'd0},p_prime[1213],s_w_1213);
AND_array_1509 AND_array_1509_c1214({a_c[294:0],1214'd0},p_prime[1214],c_w_1214);
AND_array_1509 AND_array_1509_s1214({a_s[294:0],1214'd0},p_prime[1214],s_w_1214);
AND_array_1509 AND_array_1509_c1215({a_c[293:0],1215'd0},p_prime[1215],c_w_1215);
AND_array_1509 AND_array_1509_s1215({a_s[293:0],1215'd0},p_prime[1215],s_w_1215);
AND_array_1509 AND_array_1509_c1216({a_c[292:0],1216'd0},p_prime[1216],c_w_1216);
AND_array_1509 AND_array_1509_s1216({a_s[292:0],1216'd0},p_prime[1216],s_w_1216);
AND_array_1509 AND_array_1509_c1217({a_c[291:0],1217'd0},p_prime[1217],c_w_1217);
AND_array_1509 AND_array_1509_s1217({a_s[291:0],1217'd0},p_prime[1217],s_w_1217);
AND_array_1509 AND_array_1509_c1218({a_c[290:0],1218'd0},p_prime[1218],c_w_1218);
AND_array_1509 AND_array_1509_s1218({a_s[290:0],1218'd0},p_prime[1218],s_w_1218);
AND_array_1509 AND_array_1509_c1219({a_c[289:0],1219'd0},p_prime[1219],c_w_1219);
AND_array_1509 AND_array_1509_s1219({a_s[289:0],1219'd0},p_prime[1219],s_w_1219);
AND_array_1509 AND_array_1509_c1220({a_c[288:0],1220'd0},p_prime[1220],c_w_1220);
AND_array_1509 AND_array_1509_s1220({a_s[288:0],1220'd0},p_prime[1220],s_w_1220);
AND_array_1509 AND_array_1509_c1221({a_c[287:0],1221'd0},p_prime[1221],c_w_1221);
AND_array_1509 AND_array_1509_s1221({a_s[287:0],1221'd0},p_prime[1221],s_w_1221);
AND_array_1509 AND_array_1509_c1222({a_c[286:0],1222'd0},p_prime[1222],c_w_1222);
AND_array_1509 AND_array_1509_s1222({a_s[286:0],1222'd0},p_prime[1222],s_w_1222);
AND_array_1509 AND_array_1509_c1223({a_c[285:0],1223'd0},p_prime[1223],c_w_1223);
AND_array_1509 AND_array_1509_s1223({a_s[285:0],1223'd0},p_prime[1223],s_w_1223);
AND_array_1509 AND_array_1509_c1224({a_c[284:0],1224'd0},p_prime[1224],c_w_1224);
AND_array_1509 AND_array_1509_s1224({a_s[284:0],1224'd0},p_prime[1224],s_w_1224);
AND_array_1509 AND_array_1509_c1225({a_c[283:0],1225'd0},p_prime[1225],c_w_1225);
AND_array_1509 AND_array_1509_s1225({a_s[283:0],1225'd0},p_prime[1225],s_w_1225);
AND_array_1509 AND_array_1509_c1226({a_c[282:0],1226'd0},p_prime[1226],c_w_1226);
AND_array_1509 AND_array_1509_s1226({a_s[282:0],1226'd0},p_prime[1226],s_w_1226);
AND_array_1509 AND_array_1509_c1227({a_c[281:0],1227'd0},p_prime[1227],c_w_1227);
AND_array_1509 AND_array_1509_s1227({a_s[281:0],1227'd0},p_prime[1227],s_w_1227);
AND_array_1509 AND_array_1509_c1228({a_c[280:0],1228'd0},p_prime[1228],c_w_1228);
AND_array_1509 AND_array_1509_s1228({a_s[280:0],1228'd0},p_prime[1228],s_w_1228);
AND_array_1509 AND_array_1509_c1229({a_c[279:0],1229'd0},p_prime[1229],c_w_1229);
AND_array_1509 AND_array_1509_s1229({a_s[279:0],1229'd0},p_prime[1229],s_w_1229);
AND_array_1509 AND_array_1509_c1230({a_c[278:0],1230'd0},p_prime[1230],c_w_1230);
AND_array_1509 AND_array_1509_s1230({a_s[278:0],1230'd0},p_prime[1230],s_w_1230);
AND_array_1509 AND_array_1509_c1231({a_c[277:0],1231'd0},p_prime[1231],c_w_1231);
AND_array_1509 AND_array_1509_s1231({a_s[277:0],1231'd0},p_prime[1231],s_w_1231);
AND_array_1509 AND_array_1509_c1232({a_c[276:0],1232'd0},p_prime[1232],c_w_1232);
AND_array_1509 AND_array_1509_s1232({a_s[276:0],1232'd0},p_prime[1232],s_w_1232);
AND_array_1509 AND_array_1509_c1233({a_c[275:0],1233'd0},p_prime[1233],c_w_1233);
AND_array_1509 AND_array_1509_s1233({a_s[275:0],1233'd0},p_prime[1233],s_w_1233);
AND_array_1509 AND_array_1509_c1234({a_c[274:0],1234'd0},p_prime[1234],c_w_1234);
AND_array_1509 AND_array_1509_s1234({a_s[274:0],1234'd0},p_prime[1234],s_w_1234);
AND_array_1509 AND_array_1509_c1235({a_c[273:0],1235'd0},p_prime[1235],c_w_1235);
AND_array_1509 AND_array_1509_s1235({a_s[273:0],1235'd0},p_prime[1235],s_w_1235);
AND_array_1509 AND_array_1509_c1236({a_c[272:0],1236'd0},p_prime[1236],c_w_1236);
AND_array_1509 AND_array_1509_s1236({a_s[272:0],1236'd0},p_prime[1236],s_w_1236);
AND_array_1509 AND_array_1509_c1237({a_c[271:0],1237'd0},p_prime[1237],c_w_1237);
AND_array_1509 AND_array_1509_s1237({a_s[271:0],1237'd0},p_prime[1237],s_w_1237);
AND_array_1509 AND_array_1509_c1238({a_c[270:0],1238'd0},p_prime[1238],c_w_1238);
AND_array_1509 AND_array_1509_s1238({a_s[270:0],1238'd0},p_prime[1238],s_w_1238);
AND_array_1509 AND_array_1509_c1239({a_c[269:0],1239'd0},p_prime[1239],c_w_1239);
AND_array_1509 AND_array_1509_s1239({a_s[269:0],1239'd0},p_prime[1239],s_w_1239);
AND_array_1509 AND_array_1509_c1240({a_c[268:0],1240'd0},p_prime[1240],c_w_1240);
AND_array_1509 AND_array_1509_s1240({a_s[268:0],1240'd0},p_prime[1240],s_w_1240);
AND_array_1509 AND_array_1509_c1241({a_c[267:0],1241'd0},p_prime[1241],c_w_1241);
AND_array_1509 AND_array_1509_s1241({a_s[267:0],1241'd0},p_prime[1241],s_w_1241);
AND_array_1509 AND_array_1509_c1242({a_c[266:0],1242'd0},p_prime[1242],c_w_1242);
AND_array_1509 AND_array_1509_s1242({a_s[266:0],1242'd0},p_prime[1242],s_w_1242);
AND_array_1509 AND_array_1509_c1243({a_c[265:0],1243'd0},p_prime[1243],c_w_1243);
AND_array_1509 AND_array_1509_s1243({a_s[265:0],1243'd0},p_prime[1243],s_w_1243);
AND_array_1509 AND_array_1509_c1244({a_c[264:0],1244'd0},p_prime[1244],c_w_1244);
AND_array_1509 AND_array_1509_s1244({a_s[264:0],1244'd0},p_prime[1244],s_w_1244);
AND_array_1509 AND_array_1509_c1245({a_c[263:0],1245'd0},p_prime[1245],c_w_1245);
AND_array_1509 AND_array_1509_s1245({a_s[263:0],1245'd0},p_prime[1245],s_w_1245);
AND_array_1509 AND_array_1509_c1246({a_c[262:0],1246'd0},p_prime[1246],c_w_1246);
AND_array_1509 AND_array_1509_s1246({a_s[262:0],1246'd0},p_prime[1246],s_w_1246);
AND_array_1509 AND_array_1509_c1247({a_c[261:0],1247'd0},p_prime[1247],c_w_1247);
AND_array_1509 AND_array_1509_s1247({a_s[261:0],1247'd0},p_prime[1247],s_w_1247);
AND_array_1509 AND_array_1509_c1248({a_c[260:0],1248'd0},p_prime[1248],c_w_1248);
AND_array_1509 AND_array_1509_s1248({a_s[260:0],1248'd0},p_prime[1248],s_w_1248);
AND_array_1509 AND_array_1509_c1249({a_c[259:0],1249'd0},p_prime[1249],c_w_1249);
AND_array_1509 AND_array_1509_s1249({a_s[259:0],1249'd0},p_prime[1249],s_w_1249);
AND_array_1509 AND_array_1509_c1250({a_c[258:0],1250'd0},p_prime[1250],c_w_1250);
AND_array_1509 AND_array_1509_s1250({a_s[258:0],1250'd0},p_prime[1250],s_w_1250);
AND_array_1509 AND_array_1509_c1251({a_c[257:0],1251'd0},p_prime[1251],c_w_1251);
AND_array_1509 AND_array_1509_s1251({a_s[257:0],1251'd0},p_prime[1251],s_w_1251);
AND_array_1509 AND_array_1509_c1252({a_c[256:0],1252'd0},p_prime[1252],c_w_1252);
AND_array_1509 AND_array_1509_s1252({a_s[256:0],1252'd0},p_prime[1252],s_w_1252);
AND_array_1509 AND_array_1509_c1253({a_c[255:0],1253'd0},p_prime[1253],c_w_1253);
AND_array_1509 AND_array_1509_s1253({a_s[255:0],1253'd0},p_prime[1253],s_w_1253);
AND_array_1509 AND_array_1509_c1254({a_c[254:0],1254'd0},p_prime[1254],c_w_1254);
AND_array_1509 AND_array_1509_s1254({a_s[254:0],1254'd0},p_prime[1254],s_w_1254);
AND_array_1509 AND_array_1509_c1255({a_c[253:0],1255'd0},p_prime[1255],c_w_1255);
AND_array_1509 AND_array_1509_s1255({a_s[253:0],1255'd0},p_prime[1255],s_w_1255);
AND_array_1509 AND_array_1509_c1256({a_c[252:0],1256'd0},p_prime[1256],c_w_1256);
AND_array_1509 AND_array_1509_s1256({a_s[252:0],1256'd0},p_prime[1256],s_w_1256);
AND_array_1509 AND_array_1509_c1257({a_c[251:0],1257'd0},p_prime[1257],c_w_1257);
AND_array_1509 AND_array_1509_s1257({a_s[251:0],1257'd0},p_prime[1257],s_w_1257);
AND_array_1509 AND_array_1509_c1258({a_c[250:0],1258'd0},p_prime[1258],c_w_1258);
AND_array_1509 AND_array_1509_s1258({a_s[250:0],1258'd0},p_prime[1258],s_w_1258);
AND_array_1509 AND_array_1509_c1259({a_c[249:0],1259'd0},p_prime[1259],c_w_1259);
AND_array_1509 AND_array_1509_s1259({a_s[249:0],1259'd0},p_prime[1259],s_w_1259);
AND_array_1509 AND_array_1509_c1260({a_c[248:0],1260'd0},p_prime[1260],c_w_1260);
AND_array_1509 AND_array_1509_s1260({a_s[248:0],1260'd0},p_prime[1260],s_w_1260);
AND_array_1509 AND_array_1509_c1261({a_c[247:0],1261'd0},p_prime[1261],c_w_1261);
AND_array_1509 AND_array_1509_s1261({a_s[247:0],1261'd0},p_prime[1261],s_w_1261);
AND_array_1509 AND_array_1509_c1262({a_c[246:0],1262'd0},p_prime[1262],c_w_1262);
AND_array_1509 AND_array_1509_s1262({a_s[246:0],1262'd0},p_prime[1262],s_w_1262);
AND_array_1509 AND_array_1509_c1263({a_c[245:0],1263'd0},p_prime[1263],c_w_1263);
AND_array_1509 AND_array_1509_s1263({a_s[245:0],1263'd0},p_prime[1263],s_w_1263);
AND_array_1509 AND_array_1509_c1264({a_c[244:0],1264'd0},p_prime[1264],c_w_1264);
AND_array_1509 AND_array_1509_s1264({a_s[244:0],1264'd0},p_prime[1264],s_w_1264);
AND_array_1509 AND_array_1509_c1265({a_c[243:0],1265'd0},p_prime[1265],c_w_1265);
AND_array_1509 AND_array_1509_s1265({a_s[243:0],1265'd0},p_prime[1265],s_w_1265);
AND_array_1509 AND_array_1509_c1266({a_c[242:0],1266'd0},p_prime[1266],c_w_1266);
AND_array_1509 AND_array_1509_s1266({a_s[242:0],1266'd0},p_prime[1266],s_w_1266);
AND_array_1509 AND_array_1509_c1267({a_c[241:0],1267'd0},p_prime[1267],c_w_1267);
AND_array_1509 AND_array_1509_s1267({a_s[241:0],1267'd0},p_prime[1267],s_w_1267);
AND_array_1509 AND_array_1509_c1268({a_c[240:0],1268'd0},p_prime[1268],c_w_1268);
AND_array_1509 AND_array_1509_s1268({a_s[240:0],1268'd0},p_prime[1268],s_w_1268);
AND_array_1509 AND_array_1509_c1269({a_c[239:0],1269'd0},p_prime[1269],c_w_1269);
AND_array_1509 AND_array_1509_s1269({a_s[239:0],1269'd0},p_prime[1269],s_w_1269);
AND_array_1509 AND_array_1509_c1270({a_c[238:0],1270'd0},p_prime[1270],c_w_1270);
AND_array_1509 AND_array_1509_s1270({a_s[238:0],1270'd0},p_prime[1270],s_w_1270);
AND_array_1509 AND_array_1509_c1271({a_c[237:0],1271'd0},p_prime[1271],c_w_1271);
AND_array_1509 AND_array_1509_s1271({a_s[237:0],1271'd0},p_prime[1271],s_w_1271);
AND_array_1509 AND_array_1509_c1272({a_c[236:0],1272'd0},p_prime[1272],c_w_1272);
AND_array_1509 AND_array_1509_s1272({a_s[236:0],1272'd0},p_prime[1272],s_w_1272);
AND_array_1509 AND_array_1509_c1273({a_c[235:0],1273'd0},p_prime[1273],c_w_1273);
AND_array_1509 AND_array_1509_s1273({a_s[235:0],1273'd0},p_prime[1273],s_w_1273);
AND_array_1509 AND_array_1509_c1274({a_c[234:0],1274'd0},p_prime[1274],c_w_1274);
AND_array_1509 AND_array_1509_s1274({a_s[234:0],1274'd0},p_prime[1274],s_w_1274);
AND_array_1509 AND_array_1509_c1275({a_c[233:0],1275'd0},p_prime[1275],c_w_1275);
AND_array_1509 AND_array_1509_s1275({a_s[233:0],1275'd0},p_prime[1275],s_w_1275);
AND_array_1509 AND_array_1509_c1276({a_c[232:0],1276'd0},p_prime[1276],c_w_1276);
AND_array_1509 AND_array_1509_s1276({a_s[232:0],1276'd0},p_prime[1276],s_w_1276);
AND_array_1509 AND_array_1509_c1277({a_c[231:0],1277'd0},p_prime[1277],c_w_1277);
AND_array_1509 AND_array_1509_s1277({a_s[231:0],1277'd0},p_prime[1277],s_w_1277);
AND_array_1509 AND_array_1509_c1278({a_c[230:0],1278'd0},p_prime[1278],c_w_1278);
AND_array_1509 AND_array_1509_s1278({a_s[230:0],1278'd0},p_prime[1278],s_w_1278);
AND_array_1509 AND_array_1509_c1279({a_c[229:0],1279'd0},p_prime[1279],c_w_1279);
AND_array_1509 AND_array_1509_s1279({a_s[229:0],1279'd0},p_prime[1279],s_w_1279);
AND_array_1509 AND_array_1509_c1280({a_c[228:0],1280'd0},p_prime[1280],c_w_1280);
AND_array_1509 AND_array_1509_s1280({a_s[228:0],1280'd0},p_prime[1280],s_w_1280);
AND_array_1509 AND_array_1509_c1281({a_c[227:0],1281'd0},p_prime[1281],c_w_1281);
AND_array_1509 AND_array_1509_s1281({a_s[227:0],1281'd0},p_prime[1281],s_w_1281);
AND_array_1509 AND_array_1509_c1282({a_c[226:0],1282'd0},p_prime[1282],c_w_1282);
AND_array_1509 AND_array_1509_s1282({a_s[226:0],1282'd0},p_prime[1282],s_w_1282);
AND_array_1509 AND_array_1509_c1283({a_c[225:0],1283'd0},p_prime[1283],c_w_1283);
AND_array_1509 AND_array_1509_s1283({a_s[225:0],1283'd0},p_prime[1283],s_w_1283);
AND_array_1509 AND_array_1509_c1284({a_c[224:0],1284'd0},p_prime[1284],c_w_1284);
AND_array_1509 AND_array_1509_s1284({a_s[224:0],1284'd0},p_prime[1284],s_w_1284);
AND_array_1509 AND_array_1509_c1285({a_c[223:0],1285'd0},p_prime[1285],c_w_1285);
AND_array_1509 AND_array_1509_s1285({a_s[223:0],1285'd0},p_prime[1285],s_w_1285);
AND_array_1509 AND_array_1509_c1286({a_c[222:0],1286'd0},p_prime[1286],c_w_1286);
AND_array_1509 AND_array_1509_s1286({a_s[222:0],1286'd0},p_prime[1286],s_w_1286);
AND_array_1509 AND_array_1509_c1287({a_c[221:0],1287'd0},p_prime[1287],c_w_1287);
AND_array_1509 AND_array_1509_s1287({a_s[221:0],1287'd0},p_prime[1287],s_w_1287);
AND_array_1509 AND_array_1509_c1288({a_c[220:0],1288'd0},p_prime[1288],c_w_1288);
AND_array_1509 AND_array_1509_s1288({a_s[220:0],1288'd0},p_prime[1288],s_w_1288);
AND_array_1509 AND_array_1509_c1289({a_c[219:0],1289'd0},p_prime[1289],c_w_1289);
AND_array_1509 AND_array_1509_s1289({a_s[219:0],1289'd0},p_prime[1289],s_w_1289);
AND_array_1509 AND_array_1509_c1290({a_c[218:0],1290'd0},p_prime[1290],c_w_1290);
AND_array_1509 AND_array_1509_s1290({a_s[218:0],1290'd0},p_prime[1290],s_w_1290);
AND_array_1509 AND_array_1509_c1291({a_c[217:0],1291'd0},p_prime[1291],c_w_1291);
AND_array_1509 AND_array_1509_s1291({a_s[217:0],1291'd0},p_prime[1291],s_w_1291);
AND_array_1509 AND_array_1509_c1292({a_c[216:0],1292'd0},p_prime[1292],c_w_1292);
AND_array_1509 AND_array_1509_s1292({a_s[216:0],1292'd0},p_prime[1292],s_w_1292);
AND_array_1509 AND_array_1509_c1293({a_c[215:0],1293'd0},p_prime[1293],c_w_1293);
AND_array_1509 AND_array_1509_s1293({a_s[215:0],1293'd0},p_prime[1293],s_w_1293);
AND_array_1509 AND_array_1509_c1294({a_c[214:0],1294'd0},p_prime[1294],c_w_1294);
AND_array_1509 AND_array_1509_s1294({a_s[214:0],1294'd0},p_prime[1294],s_w_1294);
AND_array_1509 AND_array_1509_c1295({a_c[213:0],1295'd0},p_prime[1295],c_w_1295);
AND_array_1509 AND_array_1509_s1295({a_s[213:0],1295'd0},p_prime[1295],s_w_1295);
AND_array_1509 AND_array_1509_c1296({a_c[212:0],1296'd0},p_prime[1296],c_w_1296);
AND_array_1509 AND_array_1509_s1296({a_s[212:0],1296'd0},p_prime[1296],s_w_1296);
AND_array_1509 AND_array_1509_c1297({a_c[211:0],1297'd0},p_prime[1297],c_w_1297);
AND_array_1509 AND_array_1509_s1297({a_s[211:0],1297'd0},p_prime[1297],s_w_1297);
AND_array_1509 AND_array_1509_c1298({a_c[210:0],1298'd0},p_prime[1298],c_w_1298);
AND_array_1509 AND_array_1509_s1298({a_s[210:0],1298'd0},p_prime[1298],s_w_1298);
AND_array_1509 AND_array_1509_c1299({a_c[209:0],1299'd0},p_prime[1299],c_w_1299);
AND_array_1509 AND_array_1509_s1299({a_s[209:0],1299'd0},p_prime[1299],s_w_1299);
AND_array_1509 AND_array_1509_c1300({a_c[208:0],1300'd0},p_prime[1300],c_w_1300);
AND_array_1509 AND_array_1509_s1300({a_s[208:0],1300'd0},p_prime[1300],s_w_1300);
AND_array_1509 AND_array_1509_c1301({a_c[207:0],1301'd0},p_prime[1301],c_w_1301);
AND_array_1509 AND_array_1509_s1301({a_s[207:0],1301'd0},p_prime[1301],s_w_1301);
AND_array_1509 AND_array_1509_c1302({a_c[206:0],1302'd0},p_prime[1302],c_w_1302);
AND_array_1509 AND_array_1509_s1302({a_s[206:0],1302'd0},p_prime[1302],s_w_1302);
AND_array_1509 AND_array_1509_c1303({a_c[205:0],1303'd0},p_prime[1303],c_w_1303);
AND_array_1509 AND_array_1509_s1303({a_s[205:0],1303'd0},p_prime[1303],s_w_1303);
AND_array_1509 AND_array_1509_c1304({a_c[204:0],1304'd0},p_prime[1304],c_w_1304);
AND_array_1509 AND_array_1509_s1304({a_s[204:0],1304'd0},p_prime[1304],s_w_1304);
AND_array_1509 AND_array_1509_c1305({a_c[203:0],1305'd0},p_prime[1305],c_w_1305);
AND_array_1509 AND_array_1509_s1305({a_s[203:0],1305'd0},p_prime[1305],s_w_1305);
AND_array_1509 AND_array_1509_c1306({a_c[202:0],1306'd0},p_prime[1306],c_w_1306);
AND_array_1509 AND_array_1509_s1306({a_s[202:0],1306'd0},p_prime[1306],s_w_1306);
AND_array_1509 AND_array_1509_c1307({a_c[201:0],1307'd0},p_prime[1307],c_w_1307);
AND_array_1509 AND_array_1509_s1307({a_s[201:0],1307'd0},p_prime[1307],s_w_1307);
AND_array_1509 AND_array_1509_c1308({a_c[200:0],1308'd0},p_prime[1308],c_w_1308);
AND_array_1509 AND_array_1509_s1308({a_s[200:0],1308'd0},p_prime[1308],s_w_1308);
AND_array_1509 AND_array_1509_c1309({a_c[199:0],1309'd0},p_prime[1309],c_w_1309);
AND_array_1509 AND_array_1509_s1309({a_s[199:0],1309'd0},p_prime[1309],s_w_1309);
AND_array_1509 AND_array_1509_c1310({a_c[198:0],1310'd0},p_prime[1310],c_w_1310);
AND_array_1509 AND_array_1509_s1310({a_s[198:0],1310'd0},p_prime[1310],s_w_1310);
AND_array_1509 AND_array_1509_c1311({a_c[197:0],1311'd0},p_prime[1311],c_w_1311);
AND_array_1509 AND_array_1509_s1311({a_s[197:0],1311'd0},p_prime[1311],s_w_1311);
AND_array_1509 AND_array_1509_c1312({a_c[196:0],1312'd0},p_prime[1312],c_w_1312);
AND_array_1509 AND_array_1509_s1312({a_s[196:0],1312'd0},p_prime[1312],s_w_1312);
AND_array_1509 AND_array_1509_c1313({a_c[195:0],1313'd0},p_prime[1313],c_w_1313);
AND_array_1509 AND_array_1509_s1313({a_s[195:0],1313'd0},p_prime[1313],s_w_1313);
AND_array_1509 AND_array_1509_c1314({a_c[194:0],1314'd0},p_prime[1314],c_w_1314);
AND_array_1509 AND_array_1509_s1314({a_s[194:0],1314'd0},p_prime[1314],s_w_1314);
AND_array_1509 AND_array_1509_c1315({a_c[193:0],1315'd0},p_prime[1315],c_w_1315);
AND_array_1509 AND_array_1509_s1315({a_s[193:0],1315'd0},p_prime[1315],s_w_1315);
AND_array_1509 AND_array_1509_c1316({a_c[192:0],1316'd0},p_prime[1316],c_w_1316);
AND_array_1509 AND_array_1509_s1316({a_s[192:0],1316'd0},p_prime[1316],s_w_1316);
AND_array_1509 AND_array_1509_c1317({a_c[191:0],1317'd0},p_prime[1317],c_w_1317);
AND_array_1509 AND_array_1509_s1317({a_s[191:0],1317'd0},p_prime[1317],s_w_1317);
AND_array_1509 AND_array_1509_c1318({a_c[190:0],1318'd0},p_prime[1318],c_w_1318);
AND_array_1509 AND_array_1509_s1318({a_s[190:0],1318'd0},p_prime[1318],s_w_1318);
AND_array_1509 AND_array_1509_c1319({a_c[189:0],1319'd0},p_prime[1319],c_w_1319);
AND_array_1509 AND_array_1509_s1319({a_s[189:0],1319'd0},p_prime[1319],s_w_1319);
AND_array_1509 AND_array_1509_c1320({a_c[188:0],1320'd0},p_prime[1320],c_w_1320);
AND_array_1509 AND_array_1509_s1320({a_s[188:0],1320'd0},p_prime[1320],s_w_1320);
AND_array_1509 AND_array_1509_c1321({a_c[187:0],1321'd0},p_prime[1321],c_w_1321);
AND_array_1509 AND_array_1509_s1321({a_s[187:0],1321'd0},p_prime[1321],s_w_1321);
AND_array_1509 AND_array_1509_c1322({a_c[186:0],1322'd0},p_prime[1322],c_w_1322);
AND_array_1509 AND_array_1509_s1322({a_s[186:0],1322'd0},p_prime[1322],s_w_1322);
AND_array_1509 AND_array_1509_c1323({a_c[185:0],1323'd0},p_prime[1323],c_w_1323);
AND_array_1509 AND_array_1509_s1323({a_s[185:0],1323'd0},p_prime[1323],s_w_1323);
AND_array_1509 AND_array_1509_c1324({a_c[184:0],1324'd0},p_prime[1324],c_w_1324);
AND_array_1509 AND_array_1509_s1324({a_s[184:0],1324'd0},p_prime[1324],s_w_1324);
AND_array_1509 AND_array_1509_c1325({a_c[183:0],1325'd0},p_prime[1325],c_w_1325);
AND_array_1509 AND_array_1509_s1325({a_s[183:0],1325'd0},p_prime[1325],s_w_1325);
AND_array_1509 AND_array_1509_c1326({a_c[182:0],1326'd0},p_prime[1326],c_w_1326);
AND_array_1509 AND_array_1509_s1326({a_s[182:0],1326'd0},p_prime[1326],s_w_1326);
AND_array_1509 AND_array_1509_c1327({a_c[181:0],1327'd0},p_prime[1327],c_w_1327);
AND_array_1509 AND_array_1509_s1327({a_s[181:0],1327'd0},p_prime[1327],s_w_1327);
AND_array_1509 AND_array_1509_c1328({a_c[180:0],1328'd0},p_prime[1328],c_w_1328);
AND_array_1509 AND_array_1509_s1328({a_s[180:0],1328'd0},p_prime[1328],s_w_1328);
AND_array_1509 AND_array_1509_c1329({a_c[179:0],1329'd0},p_prime[1329],c_w_1329);
AND_array_1509 AND_array_1509_s1329({a_s[179:0],1329'd0},p_prime[1329],s_w_1329);
AND_array_1509 AND_array_1509_c1330({a_c[178:0],1330'd0},p_prime[1330],c_w_1330);
AND_array_1509 AND_array_1509_s1330({a_s[178:0],1330'd0},p_prime[1330],s_w_1330);
AND_array_1509 AND_array_1509_c1331({a_c[177:0],1331'd0},p_prime[1331],c_w_1331);
AND_array_1509 AND_array_1509_s1331({a_s[177:0],1331'd0},p_prime[1331],s_w_1331);
AND_array_1509 AND_array_1509_c1332({a_c[176:0],1332'd0},p_prime[1332],c_w_1332);
AND_array_1509 AND_array_1509_s1332({a_s[176:0],1332'd0},p_prime[1332],s_w_1332);
AND_array_1509 AND_array_1509_c1333({a_c[175:0],1333'd0},p_prime[1333],c_w_1333);
AND_array_1509 AND_array_1509_s1333({a_s[175:0],1333'd0},p_prime[1333],s_w_1333);
AND_array_1509 AND_array_1509_c1334({a_c[174:0],1334'd0},p_prime[1334],c_w_1334);
AND_array_1509 AND_array_1509_s1334({a_s[174:0],1334'd0},p_prime[1334],s_w_1334);
AND_array_1509 AND_array_1509_c1335({a_c[173:0],1335'd0},p_prime[1335],c_w_1335);
AND_array_1509 AND_array_1509_s1335({a_s[173:0],1335'd0},p_prime[1335],s_w_1335);
AND_array_1509 AND_array_1509_c1336({a_c[172:0],1336'd0},p_prime[1336],c_w_1336);
AND_array_1509 AND_array_1509_s1336({a_s[172:0],1336'd0},p_prime[1336],s_w_1336);
AND_array_1509 AND_array_1509_c1337({a_c[171:0],1337'd0},p_prime[1337],c_w_1337);
AND_array_1509 AND_array_1509_s1337({a_s[171:0],1337'd0},p_prime[1337],s_w_1337);
AND_array_1509 AND_array_1509_c1338({a_c[170:0],1338'd0},p_prime[1338],c_w_1338);
AND_array_1509 AND_array_1509_s1338({a_s[170:0],1338'd0},p_prime[1338],s_w_1338);
AND_array_1509 AND_array_1509_c1339({a_c[169:0],1339'd0},p_prime[1339],c_w_1339);
AND_array_1509 AND_array_1509_s1339({a_s[169:0],1339'd0},p_prime[1339],s_w_1339);
AND_array_1509 AND_array_1509_c1340({a_c[168:0],1340'd0},p_prime[1340],c_w_1340);
AND_array_1509 AND_array_1509_s1340({a_s[168:0],1340'd0},p_prime[1340],s_w_1340);
AND_array_1509 AND_array_1509_c1341({a_c[167:0],1341'd0},p_prime[1341],c_w_1341);
AND_array_1509 AND_array_1509_s1341({a_s[167:0],1341'd0},p_prime[1341],s_w_1341);
AND_array_1509 AND_array_1509_c1342({a_c[166:0],1342'd0},p_prime[1342],c_w_1342);
AND_array_1509 AND_array_1509_s1342({a_s[166:0],1342'd0},p_prime[1342],s_w_1342);
AND_array_1509 AND_array_1509_c1343({a_c[165:0],1343'd0},p_prime[1343],c_w_1343);
AND_array_1509 AND_array_1509_s1343({a_s[165:0],1343'd0},p_prime[1343],s_w_1343);
AND_array_1509 AND_array_1509_c1344({a_c[164:0],1344'd0},p_prime[1344],c_w_1344);
AND_array_1509 AND_array_1509_s1344({a_s[164:0],1344'd0},p_prime[1344],s_w_1344);
AND_array_1509 AND_array_1509_c1345({a_c[163:0],1345'd0},p_prime[1345],c_w_1345);
AND_array_1509 AND_array_1509_s1345({a_s[163:0],1345'd0},p_prime[1345],s_w_1345);
AND_array_1509 AND_array_1509_c1346({a_c[162:0],1346'd0},p_prime[1346],c_w_1346);
AND_array_1509 AND_array_1509_s1346({a_s[162:0],1346'd0},p_prime[1346],s_w_1346);
AND_array_1509 AND_array_1509_c1347({a_c[161:0],1347'd0},p_prime[1347],c_w_1347);
AND_array_1509 AND_array_1509_s1347({a_s[161:0],1347'd0},p_prime[1347],s_w_1347);
AND_array_1509 AND_array_1509_c1348({a_c[160:0],1348'd0},p_prime[1348],c_w_1348);
AND_array_1509 AND_array_1509_s1348({a_s[160:0],1348'd0},p_prime[1348],s_w_1348);
AND_array_1509 AND_array_1509_c1349({a_c[159:0],1349'd0},p_prime[1349],c_w_1349);
AND_array_1509 AND_array_1509_s1349({a_s[159:0],1349'd0},p_prime[1349],s_w_1349);
AND_array_1509 AND_array_1509_c1350({a_c[158:0],1350'd0},p_prime[1350],c_w_1350);
AND_array_1509 AND_array_1509_s1350({a_s[158:0],1350'd0},p_prime[1350],s_w_1350);
AND_array_1509 AND_array_1509_c1351({a_c[157:0],1351'd0},p_prime[1351],c_w_1351);
AND_array_1509 AND_array_1509_s1351({a_s[157:0],1351'd0},p_prime[1351],s_w_1351);
AND_array_1509 AND_array_1509_c1352({a_c[156:0],1352'd0},p_prime[1352],c_w_1352);
AND_array_1509 AND_array_1509_s1352({a_s[156:0],1352'd0},p_prime[1352],s_w_1352);
AND_array_1509 AND_array_1509_c1353({a_c[155:0],1353'd0},p_prime[1353],c_w_1353);
AND_array_1509 AND_array_1509_s1353({a_s[155:0],1353'd0},p_prime[1353],s_w_1353);
AND_array_1509 AND_array_1509_c1354({a_c[154:0],1354'd0},p_prime[1354],c_w_1354);
AND_array_1509 AND_array_1509_s1354({a_s[154:0],1354'd0},p_prime[1354],s_w_1354);
AND_array_1509 AND_array_1509_c1355({a_c[153:0],1355'd0},p_prime[1355],c_w_1355);
AND_array_1509 AND_array_1509_s1355({a_s[153:0],1355'd0},p_prime[1355],s_w_1355);
AND_array_1509 AND_array_1509_c1356({a_c[152:0],1356'd0},p_prime[1356],c_w_1356);
AND_array_1509 AND_array_1509_s1356({a_s[152:0],1356'd0},p_prime[1356],s_w_1356);
AND_array_1509 AND_array_1509_c1357({a_c[151:0],1357'd0},p_prime[1357],c_w_1357);
AND_array_1509 AND_array_1509_s1357({a_s[151:0],1357'd0},p_prime[1357],s_w_1357);
AND_array_1509 AND_array_1509_c1358({a_c[150:0],1358'd0},p_prime[1358],c_w_1358);
AND_array_1509 AND_array_1509_s1358({a_s[150:0],1358'd0},p_prime[1358],s_w_1358);
AND_array_1509 AND_array_1509_c1359({a_c[149:0],1359'd0},p_prime[1359],c_w_1359);
AND_array_1509 AND_array_1509_s1359({a_s[149:0],1359'd0},p_prime[1359],s_w_1359);
AND_array_1509 AND_array_1509_c1360({a_c[148:0],1360'd0},p_prime[1360],c_w_1360);
AND_array_1509 AND_array_1509_s1360({a_s[148:0],1360'd0},p_prime[1360],s_w_1360);
AND_array_1509 AND_array_1509_c1361({a_c[147:0],1361'd0},p_prime[1361],c_w_1361);
AND_array_1509 AND_array_1509_s1361({a_s[147:0],1361'd0},p_prime[1361],s_w_1361);
AND_array_1509 AND_array_1509_c1362({a_c[146:0],1362'd0},p_prime[1362],c_w_1362);
AND_array_1509 AND_array_1509_s1362({a_s[146:0],1362'd0},p_prime[1362],s_w_1362);
AND_array_1509 AND_array_1509_c1363({a_c[145:0],1363'd0},p_prime[1363],c_w_1363);
AND_array_1509 AND_array_1509_s1363({a_s[145:0],1363'd0},p_prime[1363],s_w_1363);
AND_array_1509 AND_array_1509_c1364({a_c[144:0],1364'd0},p_prime[1364],c_w_1364);
AND_array_1509 AND_array_1509_s1364({a_s[144:0],1364'd0},p_prime[1364],s_w_1364);
AND_array_1509 AND_array_1509_c1365({a_c[143:0],1365'd0},p_prime[1365],c_w_1365);
AND_array_1509 AND_array_1509_s1365({a_s[143:0],1365'd0},p_prime[1365],s_w_1365);
AND_array_1509 AND_array_1509_c1366({a_c[142:0],1366'd0},p_prime[1366],c_w_1366);
AND_array_1509 AND_array_1509_s1366({a_s[142:0],1366'd0},p_prime[1366],s_w_1366);
AND_array_1509 AND_array_1509_c1367({a_c[141:0],1367'd0},p_prime[1367],c_w_1367);
AND_array_1509 AND_array_1509_s1367({a_s[141:0],1367'd0},p_prime[1367],s_w_1367);
AND_array_1509 AND_array_1509_c1368({a_c[140:0],1368'd0},p_prime[1368],c_w_1368);
AND_array_1509 AND_array_1509_s1368({a_s[140:0],1368'd0},p_prime[1368],s_w_1368);
AND_array_1509 AND_array_1509_c1369({a_c[139:0],1369'd0},p_prime[1369],c_w_1369);
AND_array_1509 AND_array_1509_s1369({a_s[139:0],1369'd0},p_prime[1369],s_w_1369);
AND_array_1509 AND_array_1509_c1370({a_c[138:0],1370'd0},p_prime[1370],c_w_1370);
AND_array_1509 AND_array_1509_s1370({a_s[138:0],1370'd0},p_prime[1370],s_w_1370);
AND_array_1509 AND_array_1509_c1371({a_c[137:0],1371'd0},p_prime[1371],c_w_1371);
AND_array_1509 AND_array_1509_s1371({a_s[137:0],1371'd0},p_prime[1371],s_w_1371);
AND_array_1509 AND_array_1509_c1372({a_c[136:0],1372'd0},p_prime[1372],c_w_1372);
AND_array_1509 AND_array_1509_s1372({a_s[136:0],1372'd0},p_prime[1372],s_w_1372);
AND_array_1509 AND_array_1509_c1373({a_c[135:0],1373'd0},p_prime[1373],c_w_1373);
AND_array_1509 AND_array_1509_s1373({a_s[135:0],1373'd0},p_prime[1373],s_w_1373);
AND_array_1509 AND_array_1509_c1374({a_c[134:0],1374'd0},p_prime[1374],c_w_1374);
AND_array_1509 AND_array_1509_s1374({a_s[134:0],1374'd0},p_prime[1374],s_w_1374);
AND_array_1509 AND_array_1509_c1375({a_c[133:0],1375'd0},p_prime[1375],c_w_1375);
AND_array_1509 AND_array_1509_s1375({a_s[133:0],1375'd0},p_prime[1375],s_w_1375);
AND_array_1509 AND_array_1509_c1376({a_c[132:0],1376'd0},p_prime[1376],c_w_1376);
AND_array_1509 AND_array_1509_s1376({a_s[132:0],1376'd0},p_prime[1376],s_w_1376);
AND_array_1509 AND_array_1509_c1377({a_c[131:0],1377'd0},p_prime[1377],c_w_1377);
AND_array_1509 AND_array_1509_s1377({a_s[131:0],1377'd0},p_prime[1377],s_w_1377);
AND_array_1509 AND_array_1509_c1378({a_c[130:0],1378'd0},p_prime[1378],c_w_1378);
AND_array_1509 AND_array_1509_s1378({a_s[130:0],1378'd0},p_prime[1378],s_w_1378);
AND_array_1509 AND_array_1509_c1379({a_c[129:0],1379'd0},p_prime[1379],c_w_1379);
AND_array_1509 AND_array_1509_s1379({a_s[129:0],1379'd0},p_prime[1379],s_w_1379);
AND_array_1509 AND_array_1509_c1380({a_c[128:0],1380'd0},p_prime[1380],c_w_1380);
AND_array_1509 AND_array_1509_s1380({a_s[128:0],1380'd0},p_prime[1380],s_w_1380);
AND_array_1509 AND_array_1509_c1381({a_c[127:0],1381'd0},p_prime[1381],c_w_1381);
AND_array_1509 AND_array_1509_s1381({a_s[127:0],1381'd0},p_prime[1381],s_w_1381);
AND_array_1509 AND_array_1509_c1382({a_c[126:0],1382'd0},p_prime[1382],c_w_1382);
AND_array_1509 AND_array_1509_s1382({a_s[126:0],1382'd0},p_prime[1382],s_w_1382);
AND_array_1509 AND_array_1509_c1383({a_c[125:0],1383'd0},p_prime[1383],c_w_1383);
AND_array_1509 AND_array_1509_s1383({a_s[125:0],1383'd0},p_prime[1383],s_w_1383);
AND_array_1509 AND_array_1509_c1384({a_c[124:0],1384'd0},p_prime[1384],c_w_1384);
AND_array_1509 AND_array_1509_s1384({a_s[124:0],1384'd0},p_prime[1384],s_w_1384);
AND_array_1509 AND_array_1509_c1385({a_c[123:0],1385'd0},p_prime[1385],c_w_1385);
AND_array_1509 AND_array_1509_s1385({a_s[123:0],1385'd0},p_prime[1385],s_w_1385);
AND_array_1509 AND_array_1509_c1386({a_c[122:0],1386'd0},p_prime[1386],c_w_1386);
AND_array_1509 AND_array_1509_s1386({a_s[122:0],1386'd0},p_prime[1386],s_w_1386);
AND_array_1509 AND_array_1509_c1387({a_c[121:0],1387'd0},p_prime[1387],c_w_1387);
AND_array_1509 AND_array_1509_s1387({a_s[121:0],1387'd0},p_prime[1387],s_w_1387);
AND_array_1509 AND_array_1509_c1388({a_c[120:0],1388'd0},p_prime[1388],c_w_1388);
AND_array_1509 AND_array_1509_s1388({a_s[120:0],1388'd0},p_prime[1388],s_w_1388);
AND_array_1509 AND_array_1509_c1389({a_c[119:0],1389'd0},p_prime[1389],c_w_1389);
AND_array_1509 AND_array_1509_s1389({a_s[119:0],1389'd0},p_prime[1389],s_w_1389);
AND_array_1509 AND_array_1509_c1390({a_c[118:0],1390'd0},p_prime[1390],c_w_1390);
AND_array_1509 AND_array_1509_s1390({a_s[118:0],1390'd0},p_prime[1390],s_w_1390);
AND_array_1509 AND_array_1509_c1391({a_c[117:0],1391'd0},p_prime[1391],c_w_1391);
AND_array_1509 AND_array_1509_s1391({a_s[117:0],1391'd0},p_prime[1391],s_w_1391);
AND_array_1509 AND_array_1509_c1392({a_c[116:0],1392'd0},p_prime[1392],c_w_1392);
AND_array_1509 AND_array_1509_s1392({a_s[116:0],1392'd0},p_prime[1392],s_w_1392);
AND_array_1509 AND_array_1509_c1393({a_c[115:0],1393'd0},p_prime[1393],c_w_1393);
AND_array_1509 AND_array_1509_s1393({a_s[115:0],1393'd0},p_prime[1393],s_w_1393);
AND_array_1509 AND_array_1509_c1394({a_c[114:0],1394'd0},p_prime[1394],c_w_1394);
AND_array_1509 AND_array_1509_s1394({a_s[114:0],1394'd0},p_prime[1394],s_w_1394);
AND_array_1509 AND_array_1509_c1395({a_c[113:0],1395'd0},p_prime[1395],c_w_1395);
AND_array_1509 AND_array_1509_s1395({a_s[113:0],1395'd0},p_prime[1395],s_w_1395);
AND_array_1509 AND_array_1509_c1396({a_c[112:0],1396'd0},p_prime[1396],c_w_1396);
AND_array_1509 AND_array_1509_s1396({a_s[112:0],1396'd0},p_prime[1396],s_w_1396);
AND_array_1509 AND_array_1509_c1397({a_c[111:0],1397'd0},p_prime[1397],c_w_1397);
AND_array_1509 AND_array_1509_s1397({a_s[111:0],1397'd0},p_prime[1397],s_w_1397);
AND_array_1509 AND_array_1509_c1398({a_c[110:0],1398'd0},p_prime[1398],c_w_1398);
AND_array_1509 AND_array_1509_s1398({a_s[110:0],1398'd0},p_prime[1398],s_w_1398);
AND_array_1509 AND_array_1509_c1399({a_c[109:0],1399'd0},p_prime[1399],c_w_1399);
AND_array_1509 AND_array_1509_s1399({a_s[109:0],1399'd0},p_prime[1399],s_w_1399);
AND_array_1509 AND_array_1509_c1400({a_c[108:0],1400'd0},p_prime[1400],c_w_1400);
AND_array_1509 AND_array_1509_s1400({a_s[108:0],1400'd0},p_prime[1400],s_w_1400);
AND_array_1509 AND_array_1509_c1401({a_c[107:0],1401'd0},p_prime[1401],c_w_1401);
AND_array_1509 AND_array_1509_s1401({a_s[107:0],1401'd0},p_prime[1401],s_w_1401);
AND_array_1509 AND_array_1509_c1402({a_c[106:0],1402'd0},p_prime[1402],c_w_1402);
AND_array_1509 AND_array_1509_s1402({a_s[106:0],1402'd0},p_prime[1402],s_w_1402);
AND_array_1509 AND_array_1509_c1403({a_c[105:0],1403'd0},p_prime[1403],c_w_1403);
AND_array_1509 AND_array_1509_s1403({a_s[105:0],1403'd0},p_prime[1403],s_w_1403);
AND_array_1509 AND_array_1509_c1404({a_c[104:0],1404'd0},p_prime[1404],c_w_1404);
AND_array_1509 AND_array_1509_s1404({a_s[104:0],1404'd0},p_prime[1404],s_w_1404);
AND_array_1509 AND_array_1509_c1405({a_c[103:0],1405'd0},p_prime[1405],c_w_1405);
AND_array_1509 AND_array_1509_s1405({a_s[103:0],1405'd0},p_prime[1405],s_w_1405);
AND_array_1509 AND_array_1509_c1406({a_c[102:0],1406'd0},p_prime[1406],c_w_1406);
AND_array_1509 AND_array_1509_s1406({a_s[102:0],1406'd0},p_prime[1406],s_w_1406);
AND_array_1509 AND_array_1509_c1407({a_c[101:0],1407'd0},p_prime[1407],c_w_1407);
AND_array_1509 AND_array_1509_s1407({a_s[101:0],1407'd0},p_prime[1407],s_w_1407);
AND_array_1509 AND_array_1509_c1408({a_c[100:0],1408'd0},p_prime[1408],c_w_1408);
AND_array_1509 AND_array_1509_s1408({a_s[100:0],1408'd0},p_prime[1408],s_w_1408);
AND_array_1509 AND_array_1509_c1409({a_c[99:0],1409'd0},p_prime[1409],c_w_1409);
AND_array_1509 AND_array_1509_s1409({a_s[99:0],1409'd0},p_prime[1409],s_w_1409);
AND_array_1509 AND_array_1509_c1410({a_c[98:0],1410'd0},p_prime[1410],c_w_1410);
AND_array_1509 AND_array_1509_s1410({a_s[98:0],1410'd0},p_prime[1410],s_w_1410);
AND_array_1509 AND_array_1509_c1411({a_c[97:0],1411'd0},p_prime[1411],c_w_1411);
AND_array_1509 AND_array_1509_s1411({a_s[97:0],1411'd0},p_prime[1411],s_w_1411);
AND_array_1509 AND_array_1509_c1412({a_c[96:0],1412'd0},p_prime[1412],c_w_1412);
AND_array_1509 AND_array_1509_s1412({a_s[96:0],1412'd0},p_prime[1412],s_w_1412);
AND_array_1509 AND_array_1509_c1413({a_c[95:0],1413'd0},p_prime[1413],c_w_1413);
AND_array_1509 AND_array_1509_s1413({a_s[95:0],1413'd0},p_prime[1413],s_w_1413);
AND_array_1509 AND_array_1509_c1414({a_c[94:0],1414'd0},p_prime[1414],c_w_1414);
AND_array_1509 AND_array_1509_s1414({a_s[94:0],1414'd0},p_prime[1414],s_w_1414);
AND_array_1509 AND_array_1509_c1415({a_c[93:0],1415'd0},p_prime[1415],c_w_1415);
AND_array_1509 AND_array_1509_s1415({a_s[93:0],1415'd0},p_prime[1415],s_w_1415);
AND_array_1509 AND_array_1509_c1416({a_c[92:0],1416'd0},p_prime[1416],c_w_1416);
AND_array_1509 AND_array_1509_s1416({a_s[92:0],1416'd0},p_prime[1416],s_w_1416);
AND_array_1509 AND_array_1509_c1417({a_c[91:0],1417'd0},p_prime[1417],c_w_1417);
AND_array_1509 AND_array_1509_s1417({a_s[91:0],1417'd0},p_prime[1417],s_w_1417);
AND_array_1509 AND_array_1509_c1418({a_c[90:0],1418'd0},p_prime[1418],c_w_1418);
AND_array_1509 AND_array_1509_s1418({a_s[90:0],1418'd0},p_prime[1418],s_w_1418);
AND_array_1509 AND_array_1509_c1419({a_c[89:0],1419'd0},p_prime[1419],c_w_1419);
AND_array_1509 AND_array_1509_s1419({a_s[89:0],1419'd0},p_prime[1419],s_w_1419);
AND_array_1509 AND_array_1509_c1420({a_c[88:0],1420'd0},p_prime[1420],c_w_1420);
AND_array_1509 AND_array_1509_s1420({a_s[88:0],1420'd0},p_prime[1420],s_w_1420);
AND_array_1509 AND_array_1509_c1421({a_c[87:0],1421'd0},p_prime[1421],c_w_1421);
AND_array_1509 AND_array_1509_s1421({a_s[87:0],1421'd0},p_prime[1421],s_w_1421);
AND_array_1509 AND_array_1509_c1422({a_c[86:0],1422'd0},p_prime[1422],c_w_1422);
AND_array_1509 AND_array_1509_s1422({a_s[86:0],1422'd0},p_prime[1422],s_w_1422);
AND_array_1509 AND_array_1509_c1423({a_c[85:0],1423'd0},p_prime[1423],c_w_1423);
AND_array_1509 AND_array_1509_s1423({a_s[85:0],1423'd0},p_prime[1423],s_w_1423);
AND_array_1509 AND_array_1509_c1424({a_c[84:0],1424'd0},p_prime[1424],c_w_1424);
AND_array_1509 AND_array_1509_s1424({a_s[84:0],1424'd0},p_prime[1424],s_w_1424);
AND_array_1509 AND_array_1509_c1425({a_c[83:0],1425'd0},p_prime[1425],c_w_1425);
AND_array_1509 AND_array_1509_s1425({a_s[83:0],1425'd0},p_prime[1425],s_w_1425);
AND_array_1509 AND_array_1509_c1426({a_c[82:0],1426'd0},p_prime[1426],c_w_1426);
AND_array_1509 AND_array_1509_s1426({a_s[82:0],1426'd0},p_prime[1426],s_w_1426);
AND_array_1509 AND_array_1509_c1427({a_c[81:0],1427'd0},p_prime[1427],c_w_1427);
AND_array_1509 AND_array_1509_s1427({a_s[81:0],1427'd0},p_prime[1427],s_w_1427);
AND_array_1509 AND_array_1509_c1428({a_c[80:0],1428'd0},p_prime[1428],c_w_1428);
AND_array_1509 AND_array_1509_s1428({a_s[80:0],1428'd0},p_prime[1428],s_w_1428);
AND_array_1509 AND_array_1509_c1429({a_c[79:0],1429'd0},p_prime[1429],c_w_1429);
AND_array_1509 AND_array_1509_s1429({a_s[79:0],1429'd0},p_prime[1429],s_w_1429);
AND_array_1509 AND_array_1509_c1430({a_c[78:0],1430'd0},p_prime[1430],c_w_1430);
AND_array_1509 AND_array_1509_s1430({a_s[78:0],1430'd0},p_prime[1430],s_w_1430);
AND_array_1509 AND_array_1509_c1431({a_c[77:0],1431'd0},p_prime[1431],c_w_1431);
AND_array_1509 AND_array_1509_s1431({a_s[77:0],1431'd0},p_prime[1431],s_w_1431);
AND_array_1509 AND_array_1509_c1432({a_c[76:0],1432'd0},p_prime[1432],c_w_1432);
AND_array_1509 AND_array_1509_s1432({a_s[76:0],1432'd0},p_prime[1432],s_w_1432);
AND_array_1509 AND_array_1509_c1433({a_c[75:0],1433'd0},p_prime[1433],c_w_1433);
AND_array_1509 AND_array_1509_s1433({a_s[75:0],1433'd0},p_prime[1433],s_w_1433);
AND_array_1509 AND_array_1509_c1434({a_c[74:0],1434'd0},p_prime[1434],c_w_1434);
AND_array_1509 AND_array_1509_s1434({a_s[74:0],1434'd0},p_prime[1434],s_w_1434);
AND_array_1509 AND_array_1509_c1435({a_c[73:0],1435'd0},p_prime[1435],c_w_1435);
AND_array_1509 AND_array_1509_s1435({a_s[73:0],1435'd0},p_prime[1435],s_w_1435);
AND_array_1509 AND_array_1509_c1436({a_c[72:0],1436'd0},p_prime[1436],c_w_1436);
AND_array_1509 AND_array_1509_s1436({a_s[72:0],1436'd0},p_prime[1436],s_w_1436);
AND_array_1509 AND_array_1509_c1437({a_c[71:0],1437'd0},p_prime[1437],c_w_1437);
AND_array_1509 AND_array_1509_s1437({a_s[71:0],1437'd0},p_prime[1437],s_w_1437);
AND_array_1509 AND_array_1509_c1438({a_c[70:0],1438'd0},p_prime[1438],c_w_1438);
AND_array_1509 AND_array_1509_s1438({a_s[70:0],1438'd0},p_prime[1438],s_w_1438);
AND_array_1509 AND_array_1509_c1439({a_c[69:0],1439'd0},p_prime[1439],c_w_1439);
AND_array_1509 AND_array_1509_s1439({a_s[69:0],1439'd0},p_prime[1439],s_w_1439);
AND_array_1509 AND_array_1509_c1440({a_c[68:0],1440'd0},p_prime[1440],c_w_1440);
AND_array_1509 AND_array_1509_s1440({a_s[68:0],1440'd0},p_prime[1440],s_w_1440);
AND_array_1509 AND_array_1509_c1441({a_c[67:0],1441'd0},p_prime[1441],c_w_1441);
AND_array_1509 AND_array_1509_s1441({a_s[67:0],1441'd0},p_prime[1441],s_w_1441);
AND_array_1509 AND_array_1509_c1442({a_c[66:0],1442'd0},p_prime[1442],c_w_1442);
AND_array_1509 AND_array_1509_s1442({a_s[66:0],1442'd0},p_prime[1442],s_w_1442);
AND_array_1509 AND_array_1509_c1443({a_c[65:0],1443'd0},p_prime[1443],c_w_1443);
AND_array_1509 AND_array_1509_s1443({a_s[65:0],1443'd0},p_prime[1443],s_w_1443);
AND_array_1509 AND_array_1509_c1444({a_c[64:0],1444'd0},p_prime[1444],c_w_1444);
AND_array_1509 AND_array_1509_s1444({a_s[64:0],1444'd0},p_prime[1444],s_w_1444);
AND_array_1509 AND_array_1509_c1445({a_c[63:0],1445'd0},p_prime[1445],c_w_1445);
AND_array_1509 AND_array_1509_s1445({a_s[63:0],1445'd0},p_prime[1445],s_w_1445);
AND_array_1509 AND_array_1509_c1446({a_c[62:0],1446'd0},p_prime[1446],c_w_1446);
AND_array_1509 AND_array_1509_s1446({a_s[62:0],1446'd0},p_prime[1446],s_w_1446);
AND_array_1509 AND_array_1509_c1447({a_c[61:0],1447'd0},p_prime[1447],c_w_1447);
AND_array_1509 AND_array_1509_s1447({a_s[61:0],1447'd0},p_prime[1447],s_w_1447);
AND_array_1509 AND_array_1509_c1448({a_c[60:0],1448'd0},p_prime[1448],c_w_1448);
AND_array_1509 AND_array_1509_s1448({a_s[60:0],1448'd0},p_prime[1448],s_w_1448);
AND_array_1509 AND_array_1509_c1449({a_c[59:0],1449'd0},p_prime[1449],c_w_1449);
AND_array_1509 AND_array_1509_s1449({a_s[59:0],1449'd0},p_prime[1449],s_w_1449);
AND_array_1509 AND_array_1509_c1450({a_c[58:0],1450'd0},p_prime[1450],c_w_1450);
AND_array_1509 AND_array_1509_s1450({a_s[58:0],1450'd0},p_prime[1450],s_w_1450);
AND_array_1509 AND_array_1509_c1451({a_c[57:0],1451'd0},p_prime[1451],c_w_1451);
AND_array_1509 AND_array_1509_s1451({a_s[57:0],1451'd0},p_prime[1451],s_w_1451);
AND_array_1509 AND_array_1509_c1452({a_c[56:0],1452'd0},p_prime[1452],c_w_1452);
AND_array_1509 AND_array_1509_s1452({a_s[56:0],1452'd0},p_prime[1452],s_w_1452);
AND_array_1509 AND_array_1509_c1453({a_c[55:0],1453'd0},p_prime[1453],c_w_1453);
AND_array_1509 AND_array_1509_s1453({a_s[55:0],1453'd0},p_prime[1453],s_w_1453);
AND_array_1509 AND_array_1509_c1454({a_c[54:0],1454'd0},p_prime[1454],c_w_1454);
AND_array_1509 AND_array_1509_s1454({a_s[54:0],1454'd0},p_prime[1454],s_w_1454);
AND_array_1509 AND_array_1509_c1455({a_c[53:0],1455'd0},p_prime[1455],c_w_1455);
AND_array_1509 AND_array_1509_s1455({a_s[53:0],1455'd0},p_prime[1455],s_w_1455);
AND_array_1509 AND_array_1509_c1456({a_c[52:0],1456'd0},p_prime[1456],c_w_1456);
AND_array_1509 AND_array_1509_s1456({a_s[52:0],1456'd0},p_prime[1456],s_w_1456);
AND_array_1509 AND_array_1509_c1457({a_c[51:0],1457'd0},p_prime[1457],c_w_1457);
AND_array_1509 AND_array_1509_s1457({a_s[51:0],1457'd0},p_prime[1457],s_w_1457);
AND_array_1509 AND_array_1509_c1458({a_c[50:0],1458'd0},p_prime[1458],c_w_1458);
AND_array_1509 AND_array_1509_s1458({a_s[50:0],1458'd0},p_prime[1458],s_w_1458);
AND_array_1509 AND_array_1509_c1459({a_c[49:0],1459'd0},p_prime[1459],c_w_1459);
AND_array_1509 AND_array_1509_s1459({a_s[49:0],1459'd0},p_prime[1459],s_w_1459);
AND_array_1509 AND_array_1509_c1460({a_c[48:0],1460'd0},p_prime[1460],c_w_1460);
AND_array_1509 AND_array_1509_s1460({a_s[48:0],1460'd0},p_prime[1460],s_w_1460);
AND_array_1509 AND_array_1509_c1461({a_c[47:0],1461'd0},p_prime[1461],c_w_1461);
AND_array_1509 AND_array_1509_s1461({a_s[47:0],1461'd0},p_prime[1461],s_w_1461);
AND_array_1509 AND_array_1509_c1462({a_c[46:0],1462'd0},p_prime[1462],c_w_1462);
AND_array_1509 AND_array_1509_s1462({a_s[46:0],1462'd0},p_prime[1462],s_w_1462);
AND_array_1509 AND_array_1509_c1463({a_c[45:0],1463'd0},p_prime[1463],c_w_1463);
AND_array_1509 AND_array_1509_s1463({a_s[45:0],1463'd0},p_prime[1463],s_w_1463);
AND_array_1509 AND_array_1509_c1464({a_c[44:0],1464'd0},p_prime[1464],c_w_1464);
AND_array_1509 AND_array_1509_s1464({a_s[44:0],1464'd0},p_prime[1464],s_w_1464);
AND_array_1509 AND_array_1509_c1465({a_c[43:0],1465'd0},p_prime[1465],c_w_1465);
AND_array_1509 AND_array_1509_s1465({a_s[43:0],1465'd0},p_prime[1465],s_w_1465);
AND_array_1509 AND_array_1509_c1466({a_c[42:0],1466'd0},p_prime[1466],c_w_1466);
AND_array_1509 AND_array_1509_s1466({a_s[42:0],1466'd0},p_prime[1466],s_w_1466);
AND_array_1509 AND_array_1509_c1467({a_c[41:0],1467'd0},p_prime[1467],c_w_1467);
AND_array_1509 AND_array_1509_s1467({a_s[41:0],1467'd0},p_prime[1467],s_w_1467);
AND_array_1509 AND_array_1509_c1468({a_c[40:0],1468'd0},p_prime[1468],c_w_1468);
AND_array_1509 AND_array_1509_s1468({a_s[40:0],1468'd0},p_prime[1468],s_w_1468);
AND_array_1509 AND_array_1509_c1469({a_c[39:0],1469'd0},p_prime[1469],c_w_1469);
AND_array_1509 AND_array_1509_s1469({a_s[39:0],1469'd0},p_prime[1469],s_w_1469);
AND_array_1509 AND_array_1509_c1470({a_c[38:0],1470'd0},p_prime[1470],c_w_1470);
AND_array_1509 AND_array_1509_s1470({a_s[38:0],1470'd0},p_prime[1470],s_w_1470);
AND_array_1509 AND_array_1509_c1471({a_c[37:0],1471'd0},p_prime[1471],c_w_1471);
AND_array_1509 AND_array_1509_s1471({a_s[37:0],1471'd0},p_prime[1471],s_w_1471);
AND_array_1509 AND_array_1509_c1472({a_c[36:0],1472'd0},p_prime[1472],c_w_1472);
AND_array_1509 AND_array_1509_s1472({a_s[36:0],1472'd0},p_prime[1472],s_w_1472);
AND_array_1509 AND_array_1509_c1473({a_c[35:0],1473'd0},p_prime[1473],c_w_1473);
AND_array_1509 AND_array_1509_s1473({a_s[35:0],1473'd0},p_prime[1473],s_w_1473);
AND_array_1509 AND_array_1509_c1474({a_c[34:0],1474'd0},p_prime[1474],c_w_1474);
AND_array_1509 AND_array_1509_s1474({a_s[34:0],1474'd0},p_prime[1474],s_w_1474);
AND_array_1509 AND_array_1509_c1475({a_c[33:0],1475'd0},p_prime[1475],c_w_1475);
AND_array_1509 AND_array_1509_s1475({a_s[33:0],1475'd0},p_prime[1475],s_w_1475);
AND_array_1509 AND_array_1509_c1476({a_c[32:0],1476'd0},p_prime[1476],c_w_1476);
AND_array_1509 AND_array_1509_s1476({a_s[32:0],1476'd0},p_prime[1476],s_w_1476);
AND_array_1509 AND_array_1509_c1477({a_c[31:0],1477'd0},p_prime[1477],c_w_1477);
AND_array_1509 AND_array_1509_s1477({a_s[31:0],1477'd0},p_prime[1477],s_w_1477);
AND_array_1509 AND_array_1509_c1478({a_c[30:0],1478'd0},p_prime[1478],c_w_1478);
AND_array_1509 AND_array_1509_s1478({a_s[30:0],1478'd0},p_prime[1478],s_w_1478);
AND_array_1509 AND_array_1509_c1479({a_c[29:0],1479'd0},p_prime[1479],c_w_1479);
AND_array_1509 AND_array_1509_s1479({a_s[29:0],1479'd0},p_prime[1479],s_w_1479);
AND_array_1509 AND_array_1509_c1480({a_c[28:0],1480'd0},p_prime[1480],c_w_1480);
AND_array_1509 AND_array_1509_s1480({a_s[28:0],1480'd0},p_prime[1480],s_w_1480);
AND_array_1509 AND_array_1509_c1481({a_c[27:0],1481'd0},p_prime[1481],c_w_1481);
AND_array_1509 AND_array_1509_s1481({a_s[27:0],1481'd0},p_prime[1481],s_w_1481);
AND_array_1509 AND_array_1509_c1482({a_c[26:0],1482'd0},p_prime[1482],c_w_1482);
AND_array_1509 AND_array_1509_s1482({a_s[26:0],1482'd0},p_prime[1482],s_w_1482);
AND_array_1509 AND_array_1509_c1483({a_c[25:0],1483'd0},p_prime[1483],c_w_1483);
AND_array_1509 AND_array_1509_s1483({a_s[25:0],1483'd0},p_prime[1483],s_w_1483);
AND_array_1509 AND_array_1509_c1484({a_c[24:0],1484'd0},p_prime[1484],c_w_1484);
AND_array_1509 AND_array_1509_s1484({a_s[24:0],1484'd0},p_prime[1484],s_w_1484);
AND_array_1509 AND_array_1509_c1485({a_c[23:0],1485'd0},p_prime[1485],c_w_1485);
AND_array_1509 AND_array_1509_s1485({a_s[23:0],1485'd0},p_prime[1485],s_w_1485);
AND_array_1509 AND_array_1509_c1486({a_c[22:0],1486'd0},p_prime[1486],c_w_1486);
AND_array_1509 AND_array_1509_s1486({a_s[22:0],1486'd0},p_prime[1486],s_w_1486);
AND_array_1509 AND_array_1509_c1487({a_c[21:0],1487'd0},p_prime[1487],c_w_1487);
AND_array_1509 AND_array_1509_s1487({a_s[21:0],1487'd0},p_prime[1487],s_w_1487);
AND_array_1509 AND_array_1509_c1488({a_c[20:0],1488'd0},p_prime[1488],c_w_1488);
AND_array_1509 AND_array_1509_s1488({a_s[20:0],1488'd0},p_prime[1488],s_w_1488);
AND_array_1509 AND_array_1509_c1489({a_c[19:0],1489'd0},p_prime[1489],c_w_1489);
AND_array_1509 AND_array_1509_s1489({a_s[19:0],1489'd0},p_prime[1489],s_w_1489);
AND_array_1509 AND_array_1509_c1490({a_c[18:0],1490'd0},p_prime[1490],c_w_1490);
AND_array_1509 AND_array_1509_s1490({a_s[18:0],1490'd0},p_prime[1490],s_w_1490);
AND_array_1509 AND_array_1509_c1491({a_c[17:0],1491'd0},p_prime[1491],c_w_1491);
AND_array_1509 AND_array_1509_s1491({a_s[17:0],1491'd0},p_prime[1491],s_w_1491);
AND_array_1509 AND_array_1509_c1492({a_c[16:0],1492'd0},p_prime[1492],c_w_1492);
AND_array_1509 AND_array_1509_s1492({a_s[16:0],1492'd0},p_prime[1492],s_w_1492);
AND_array_1509 AND_array_1509_c1493({a_c[15:0],1493'd0},p_prime[1493],c_w_1493);
AND_array_1509 AND_array_1509_s1493({a_s[15:0],1493'd0},p_prime[1493],s_w_1493);
AND_array_1509 AND_array_1509_c1494({a_c[14:0],1494'd0},p_prime[1494],c_w_1494);
AND_array_1509 AND_array_1509_s1494({a_s[14:0],1494'd0},p_prime[1494],s_w_1494);
AND_array_1509 AND_array_1509_c1495({a_c[13:0],1495'd0},p_prime[1495],c_w_1495);
AND_array_1509 AND_array_1509_s1495({a_s[13:0],1495'd0},p_prime[1495],s_w_1495);
AND_array_1509 AND_array_1509_c1496({a_c[12:0],1496'd0},p_prime[1496],c_w_1496);
AND_array_1509 AND_array_1509_s1496({a_s[12:0],1496'd0},p_prime[1496],s_w_1496);
AND_array_1509 AND_array_1509_c1497({a_c[11:0],1497'd0},p_prime[1497],c_w_1497);
AND_array_1509 AND_array_1509_s1497({a_s[11:0],1497'd0},p_prime[1497],s_w_1497);
AND_array_1509 AND_array_1509_c1498({a_c[10:0],1498'd0},p_prime[1498],c_w_1498);
AND_array_1509 AND_array_1509_s1498({a_s[10:0],1498'd0},p_prime[1498],s_w_1498);
AND_array_1509 AND_array_1509_c1499({a_c[9:0],1499'd0},p_prime[1499],c_w_1499);
AND_array_1509 AND_array_1509_s1499({a_s[9:0],1499'd0},p_prime[1499],s_w_1499);
AND_array_1509 AND_array_1509_c1500({a_c[8:0],1500'd0},p_prime[1500],c_w_1500);
AND_array_1509 AND_array_1509_s1500({a_s[8:0],1500'd0},p_prime[1500],s_w_1500);
AND_array_1509 AND_array_1509_c1501({a_c[7:0],1501'd0},p_prime[1501],c_w_1501);
AND_array_1509 AND_array_1509_s1501({a_s[7:0],1501'd0},p_prime[1501],s_w_1501);
AND_array_1509 AND_array_1509_c1502({a_c[6:0],1502'd0},p_prime[1502],c_w_1502);
AND_array_1509 AND_array_1509_s1502({a_s[6:0],1502'd0},p_prime[1502],s_w_1502);
AND_array_1509 AND_array_1509_c1503({a_c[5:0],1503'd0},p_prime[1503],c_w_1503);
AND_array_1509 AND_array_1509_s1503({a_s[5:0],1503'd0},p_prime[1503],s_w_1503);
AND_array_1509 AND_array_1509_c1504({a_c[4:0],1504'd0},p_prime[1504],c_w_1504);
AND_array_1509 AND_array_1509_s1504({a_s[4:0],1504'd0},p_prime[1504],s_w_1504);
AND_array_1509 AND_array_1509_c1505({a_c[3:0],1505'd0},p_prime[1505],c_w_1505);
AND_array_1509 AND_array_1509_s1505({a_s[3:0],1505'd0},p_prime[1505],s_w_1505);
AND_array_1509 AND_array_1509_c1506({a_c[2:0],1506'd0},p_prime[1506],c_w_1506);
AND_array_1509 AND_array_1509_s1506({a_s[2:0],1506'd0},p_prime[1506],s_w_1506);
AND_array_1509 AND_array_1509_c1507({a_c[1:0],1507'd0},p_prime[1507],c_w_1507);
AND_array_1509 AND_array_1509_s1507({a_s[1:0],1507'd0},p_prime[1507],s_w_1507);
AND_array_1509 AND_array_1509_c1508({a_c[0:0],1508'd0},p_prime[1508],c_w_1508);
AND_array_1509 AND_array_1509_s1508({a_s[0:0],1508'd0},p_prime[1508],s_w_1508);
    
assign b_c[1508:0] = c_w_0;assign b_s[1508:0] = s_w_0;
assign b_c[3017:1509] = c_w_1;assign b_s[3017:1509] = s_w_1;
assign b_c[4526:3018] = c_w_2;assign b_s[4526:3018] = s_w_2;
assign b_c[6035:4527] = c_w_3;assign b_s[6035:4527] = s_w_3;
assign b_c[7544:6036] = c_w_4;assign b_s[7544:6036] = s_w_4;
assign b_c[9053:7545] = c_w_5;assign b_s[9053:7545] = s_w_5;
assign b_c[10562:9054] = c_w_6;assign b_s[10562:9054] = s_w_6;
assign b_c[12071:10563] = c_w_7;assign b_s[12071:10563] = s_w_7;
assign b_c[13580:12072] = c_w_8;assign b_s[13580:12072] = s_w_8;
assign b_c[15089:13581] = c_w_9;assign b_s[15089:13581] = s_w_9;
assign b_c[16598:15090] = c_w_10;assign b_s[16598:15090] = s_w_10;
assign b_c[18107:16599] = c_w_11;assign b_s[18107:16599] = s_w_11;
assign b_c[19616:18108] = c_w_12;assign b_s[19616:18108] = s_w_12;
assign b_c[21125:19617] = c_w_13;assign b_s[21125:19617] = s_w_13;
assign b_c[22634:21126] = c_w_14;assign b_s[22634:21126] = s_w_14;
assign b_c[24143:22635] = c_w_15;assign b_s[24143:22635] = s_w_15;
assign b_c[25652:24144] = c_w_16;assign b_s[25652:24144] = s_w_16;
assign b_c[27161:25653] = c_w_17;assign b_s[27161:25653] = s_w_17;
assign b_c[28670:27162] = c_w_18;assign b_s[28670:27162] = s_w_18;
assign b_c[30179:28671] = c_w_19;assign b_s[30179:28671] = s_w_19;
assign b_c[31688:30180] = c_w_20;assign b_s[31688:30180] = s_w_20;
assign b_c[33197:31689] = c_w_21;assign b_s[33197:31689] = s_w_21;
assign b_c[34706:33198] = c_w_22;assign b_s[34706:33198] = s_w_22;
assign b_c[36215:34707] = c_w_23;assign b_s[36215:34707] = s_w_23;
assign b_c[37724:36216] = c_w_24;assign b_s[37724:36216] = s_w_24;
assign b_c[39233:37725] = c_w_25;assign b_s[39233:37725] = s_w_25;
assign b_c[40742:39234] = c_w_26;assign b_s[40742:39234] = s_w_26;
assign b_c[42251:40743] = c_w_27;assign b_s[42251:40743] = s_w_27;
assign b_c[43760:42252] = c_w_28;assign b_s[43760:42252] = s_w_28;
assign b_c[45269:43761] = c_w_29;assign b_s[45269:43761] = s_w_29;
assign b_c[46778:45270] = c_w_30;assign b_s[46778:45270] = s_w_30;
assign b_c[48287:46779] = c_w_31;assign b_s[48287:46779] = s_w_31;
assign b_c[49796:48288] = c_w_32;assign b_s[49796:48288] = s_w_32;
assign b_c[51305:49797] = c_w_33;assign b_s[51305:49797] = s_w_33;
assign b_c[52814:51306] = c_w_34;assign b_s[52814:51306] = s_w_34;
assign b_c[54323:52815] = c_w_35;assign b_s[54323:52815] = s_w_35;
assign b_c[55832:54324] = c_w_36;assign b_s[55832:54324] = s_w_36;
assign b_c[57341:55833] = c_w_37;assign b_s[57341:55833] = s_w_37;
assign b_c[58850:57342] = c_w_38;assign b_s[58850:57342] = s_w_38;
assign b_c[60359:58851] = c_w_39;assign b_s[60359:58851] = s_w_39;
assign b_c[61868:60360] = c_w_40;assign b_s[61868:60360] = s_w_40;
assign b_c[63377:61869] = c_w_41;assign b_s[63377:61869] = s_w_41;
assign b_c[64886:63378] = c_w_42;assign b_s[64886:63378] = s_w_42;
assign b_c[66395:64887] = c_w_43;assign b_s[66395:64887] = s_w_43;
assign b_c[67904:66396] = c_w_44;assign b_s[67904:66396] = s_w_44;
assign b_c[69413:67905] = c_w_45;assign b_s[69413:67905] = s_w_45;
assign b_c[70922:69414] = c_w_46;assign b_s[70922:69414] = s_w_46;
assign b_c[72431:70923] = c_w_47;assign b_s[72431:70923] = s_w_47;
assign b_c[73940:72432] = c_w_48;assign b_s[73940:72432] = s_w_48;
assign b_c[75449:73941] = c_w_49;assign b_s[75449:73941] = s_w_49;
assign b_c[76958:75450] = c_w_50;assign b_s[76958:75450] = s_w_50;
assign b_c[78467:76959] = c_w_51;assign b_s[78467:76959] = s_w_51;
assign b_c[79976:78468] = c_w_52;assign b_s[79976:78468] = s_w_52;
assign b_c[81485:79977] = c_w_53;assign b_s[81485:79977] = s_w_53;
assign b_c[82994:81486] = c_w_54;assign b_s[82994:81486] = s_w_54;
assign b_c[84503:82995] = c_w_55;assign b_s[84503:82995] = s_w_55;
assign b_c[86012:84504] = c_w_56;assign b_s[86012:84504] = s_w_56;
assign b_c[87521:86013] = c_w_57;assign b_s[87521:86013] = s_w_57;
assign b_c[89030:87522] = c_w_58;assign b_s[89030:87522] = s_w_58;
assign b_c[90539:89031] = c_w_59;assign b_s[90539:89031] = s_w_59;
assign b_c[92048:90540] = c_w_60;assign b_s[92048:90540] = s_w_60;
assign b_c[93557:92049] = c_w_61;assign b_s[93557:92049] = s_w_61;
assign b_c[95066:93558] = c_w_62;assign b_s[95066:93558] = s_w_62;
assign b_c[96575:95067] = c_w_63;assign b_s[96575:95067] = s_w_63;
assign b_c[98084:96576] = c_w_64;assign b_s[98084:96576] = s_w_64;
assign b_c[99593:98085] = c_w_65;assign b_s[99593:98085] = s_w_65;
assign b_c[101102:99594] = c_w_66;assign b_s[101102:99594] = s_w_66;
assign b_c[102611:101103] = c_w_67;assign b_s[102611:101103] = s_w_67;
assign b_c[104120:102612] = c_w_68;assign b_s[104120:102612] = s_w_68;
assign b_c[105629:104121] = c_w_69;assign b_s[105629:104121] = s_w_69;
assign b_c[107138:105630] = c_w_70;assign b_s[107138:105630] = s_w_70;
assign b_c[108647:107139] = c_w_71;assign b_s[108647:107139] = s_w_71;
assign b_c[110156:108648] = c_w_72;assign b_s[110156:108648] = s_w_72;
assign b_c[111665:110157] = c_w_73;assign b_s[111665:110157] = s_w_73;
assign b_c[113174:111666] = c_w_74;assign b_s[113174:111666] = s_w_74;
assign b_c[114683:113175] = c_w_75;assign b_s[114683:113175] = s_w_75;
assign b_c[116192:114684] = c_w_76;assign b_s[116192:114684] = s_w_76;
assign b_c[117701:116193] = c_w_77;assign b_s[117701:116193] = s_w_77;
assign b_c[119210:117702] = c_w_78;assign b_s[119210:117702] = s_w_78;
assign b_c[120719:119211] = c_w_79;assign b_s[120719:119211] = s_w_79;
assign b_c[122228:120720] = c_w_80;assign b_s[122228:120720] = s_w_80;
assign b_c[123737:122229] = c_w_81;assign b_s[123737:122229] = s_w_81;
assign b_c[125246:123738] = c_w_82;assign b_s[125246:123738] = s_w_82;
assign b_c[126755:125247] = c_w_83;assign b_s[126755:125247] = s_w_83;
assign b_c[128264:126756] = c_w_84;assign b_s[128264:126756] = s_w_84;
assign b_c[129773:128265] = c_w_85;assign b_s[129773:128265] = s_w_85;
assign b_c[131282:129774] = c_w_86;assign b_s[131282:129774] = s_w_86;
assign b_c[132791:131283] = c_w_87;assign b_s[132791:131283] = s_w_87;
assign b_c[134300:132792] = c_w_88;assign b_s[134300:132792] = s_w_88;
assign b_c[135809:134301] = c_w_89;assign b_s[135809:134301] = s_w_89;
assign b_c[137318:135810] = c_w_90;assign b_s[137318:135810] = s_w_90;
assign b_c[138827:137319] = c_w_91;assign b_s[138827:137319] = s_w_91;
assign b_c[140336:138828] = c_w_92;assign b_s[140336:138828] = s_w_92;
assign b_c[141845:140337] = c_w_93;assign b_s[141845:140337] = s_w_93;
assign b_c[143354:141846] = c_w_94;assign b_s[143354:141846] = s_w_94;
assign b_c[144863:143355] = c_w_95;assign b_s[144863:143355] = s_w_95;
assign b_c[146372:144864] = c_w_96;assign b_s[146372:144864] = s_w_96;
assign b_c[147881:146373] = c_w_97;assign b_s[147881:146373] = s_w_97;
assign b_c[149390:147882] = c_w_98;assign b_s[149390:147882] = s_w_98;
assign b_c[150899:149391] = c_w_99;assign b_s[150899:149391] = s_w_99;
assign b_c[152408:150900] = c_w_100;assign b_s[152408:150900] = s_w_100;
assign b_c[153917:152409] = c_w_101;assign b_s[153917:152409] = s_w_101;
assign b_c[155426:153918] = c_w_102;assign b_s[155426:153918] = s_w_102;
assign b_c[156935:155427] = c_w_103;assign b_s[156935:155427] = s_w_103;
assign b_c[158444:156936] = c_w_104;assign b_s[158444:156936] = s_w_104;
assign b_c[159953:158445] = c_w_105;assign b_s[159953:158445] = s_w_105;
assign b_c[161462:159954] = c_w_106;assign b_s[161462:159954] = s_w_106;
assign b_c[162971:161463] = c_w_107;assign b_s[162971:161463] = s_w_107;
assign b_c[164480:162972] = c_w_108;assign b_s[164480:162972] = s_w_108;
assign b_c[165989:164481] = c_w_109;assign b_s[165989:164481] = s_w_109;
assign b_c[167498:165990] = c_w_110;assign b_s[167498:165990] = s_w_110;
assign b_c[169007:167499] = c_w_111;assign b_s[169007:167499] = s_w_111;
assign b_c[170516:169008] = c_w_112;assign b_s[170516:169008] = s_w_112;
assign b_c[172025:170517] = c_w_113;assign b_s[172025:170517] = s_w_113;
assign b_c[173534:172026] = c_w_114;assign b_s[173534:172026] = s_w_114;
assign b_c[175043:173535] = c_w_115;assign b_s[175043:173535] = s_w_115;
assign b_c[176552:175044] = c_w_116;assign b_s[176552:175044] = s_w_116;
assign b_c[178061:176553] = c_w_117;assign b_s[178061:176553] = s_w_117;
assign b_c[179570:178062] = c_w_118;assign b_s[179570:178062] = s_w_118;
assign b_c[181079:179571] = c_w_119;assign b_s[181079:179571] = s_w_119;
assign b_c[182588:181080] = c_w_120;assign b_s[182588:181080] = s_w_120;
assign b_c[184097:182589] = c_w_121;assign b_s[184097:182589] = s_w_121;
assign b_c[185606:184098] = c_w_122;assign b_s[185606:184098] = s_w_122;
assign b_c[187115:185607] = c_w_123;assign b_s[187115:185607] = s_w_123;
assign b_c[188624:187116] = c_w_124;assign b_s[188624:187116] = s_w_124;
assign b_c[190133:188625] = c_w_125;assign b_s[190133:188625] = s_w_125;
assign b_c[191642:190134] = c_w_126;assign b_s[191642:190134] = s_w_126;
assign b_c[193151:191643] = c_w_127;assign b_s[193151:191643] = s_w_127;
assign b_c[194660:193152] = c_w_128;assign b_s[194660:193152] = s_w_128;
assign b_c[196169:194661] = c_w_129;assign b_s[196169:194661] = s_w_129;
assign b_c[197678:196170] = c_w_130;assign b_s[197678:196170] = s_w_130;
assign b_c[199187:197679] = c_w_131;assign b_s[199187:197679] = s_w_131;
assign b_c[200696:199188] = c_w_132;assign b_s[200696:199188] = s_w_132;
assign b_c[202205:200697] = c_w_133;assign b_s[202205:200697] = s_w_133;
assign b_c[203714:202206] = c_w_134;assign b_s[203714:202206] = s_w_134;
assign b_c[205223:203715] = c_w_135;assign b_s[205223:203715] = s_w_135;
assign b_c[206732:205224] = c_w_136;assign b_s[206732:205224] = s_w_136;
assign b_c[208241:206733] = c_w_137;assign b_s[208241:206733] = s_w_137;
assign b_c[209750:208242] = c_w_138;assign b_s[209750:208242] = s_w_138;
assign b_c[211259:209751] = c_w_139;assign b_s[211259:209751] = s_w_139;
assign b_c[212768:211260] = c_w_140;assign b_s[212768:211260] = s_w_140;
assign b_c[214277:212769] = c_w_141;assign b_s[214277:212769] = s_w_141;
assign b_c[215786:214278] = c_w_142;assign b_s[215786:214278] = s_w_142;
assign b_c[217295:215787] = c_w_143;assign b_s[217295:215787] = s_w_143;
assign b_c[218804:217296] = c_w_144;assign b_s[218804:217296] = s_w_144;
assign b_c[220313:218805] = c_w_145;assign b_s[220313:218805] = s_w_145;
assign b_c[221822:220314] = c_w_146;assign b_s[221822:220314] = s_w_146;
assign b_c[223331:221823] = c_w_147;assign b_s[223331:221823] = s_w_147;
assign b_c[224840:223332] = c_w_148;assign b_s[224840:223332] = s_w_148;
assign b_c[226349:224841] = c_w_149;assign b_s[226349:224841] = s_w_149;
assign b_c[227858:226350] = c_w_150;assign b_s[227858:226350] = s_w_150;
assign b_c[229367:227859] = c_w_151;assign b_s[229367:227859] = s_w_151;
assign b_c[230876:229368] = c_w_152;assign b_s[230876:229368] = s_w_152;
assign b_c[232385:230877] = c_w_153;assign b_s[232385:230877] = s_w_153;
assign b_c[233894:232386] = c_w_154;assign b_s[233894:232386] = s_w_154;
assign b_c[235403:233895] = c_w_155;assign b_s[235403:233895] = s_w_155;
assign b_c[236912:235404] = c_w_156;assign b_s[236912:235404] = s_w_156;
assign b_c[238421:236913] = c_w_157;assign b_s[238421:236913] = s_w_157;
assign b_c[239930:238422] = c_w_158;assign b_s[239930:238422] = s_w_158;
assign b_c[241439:239931] = c_w_159;assign b_s[241439:239931] = s_w_159;
assign b_c[242948:241440] = c_w_160;assign b_s[242948:241440] = s_w_160;
assign b_c[244457:242949] = c_w_161;assign b_s[244457:242949] = s_w_161;
assign b_c[245966:244458] = c_w_162;assign b_s[245966:244458] = s_w_162;
assign b_c[247475:245967] = c_w_163;assign b_s[247475:245967] = s_w_163;
assign b_c[248984:247476] = c_w_164;assign b_s[248984:247476] = s_w_164;
assign b_c[250493:248985] = c_w_165;assign b_s[250493:248985] = s_w_165;
assign b_c[252002:250494] = c_w_166;assign b_s[252002:250494] = s_w_166;
assign b_c[253511:252003] = c_w_167;assign b_s[253511:252003] = s_w_167;
assign b_c[255020:253512] = c_w_168;assign b_s[255020:253512] = s_w_168;
assign b_c[256529:255021] = c_w_169;assign b_s[256529:255021] = s_w_169;
assign b_c[258038:256530] = c_w_170;assign b_s[258038:256530] = s_w_170;
assign b_c[259547:258039] = c_w_171;assign b_s[259547:258039] = s_w_171;
assign b_c[261056:259548] = c_w_172;assign b_s[261056:259548] = s_w_172;
assign b_c[262565:261057] = c_w_173;assign b_s[262565:261057] = s_w_173;
assign b_c[264074:262566] = c_w_174;assign b_s[264074:262566] = s_w_174;
assign b_c[265583:264075] = c_w_175;assign b_s[265583:264075] = s_w_175;
assign b_c[267092:265584] = c_w_176;assign b_s[267092:265584] = s_w_176;
assign b_c[268601:267093] = c_w_177;assign b_s[268601:267093] = s_w_177;
assign b_c[270110:268602] = c_w_178;assign b_s[270110:268602] = s_w_178;
assign b_c[271619:270111] = c_w_179;assign b_s[271619:270111] = s_w_179;
assign b_c[273128:271620] = c_w_180;assign b_s[273128:271620] = s_w_180;
assign b_c[274637:273129] = c_w_181;assign b_s[274637:273129] = s_w_181;
assign b_c[276146:274638] = c_w_182;assign b_s[276146:274638] = s_w_182;
assign b_c[277655:276147] = c_w_183;assign b_s[277655:276147] = s_w_183;
assign b_c[279164:277656] = c_w_184;assign b_s[279164:277656] = s_w_184;
assign b_c[280673:279165] = c_w_185;assign b_s[280673:279165] = s_w_185;
assign b_c[282182:280674] = c_w_186;assign b_s[282182:280674] = s_w_186;
assign b_c[283691:282183] = c_w_187;assign b_s[283691:282183] = s_w_187;
assign b_c[285200:283692] = c_w_188;assign b_s[285200:283692] = s_w_188;
assign b_c[286709:285201] = c_w_189;assign b_s[286709:285201] = s_w_189;
assign b_c[288218:286710] = c_w_190;assign b_s[288218:286710] = s_w_190;
assign b_c[289727:288219] = c_w_191;assign b_s[289727:288219] = s_w_191;
assign b_c[291236:289728] = c_w_192;assign b_s[291236:289728] = s_w_192;
assign b_c[292745:291237] = c_w_193;assign b_s[292745:291237] = s_w_193;
assign b_c[294254:292746] = c_w_194;assign b_s[294254:292746] = s_w_194;
assign b_c[295763:294255] = c_w_195;assign b_s[295763:294255] = s_w_195;
assign b_c[297272:295764] = c_w_196;assign b_s[297272:295764] = s_w_196;
assign b_c[298781:297273] = c_w_197;assign b_s[298781:297273] = s_w_197;
assign b_c[300290:298782] = c_w_198;assign b_s[300290:298782] = s_w_198;
assign b_c[301799:300291] = c_w_199;assign b_s[301799:300291] = s_w_199;
assign b_c[303308:301800] = c_w_200;assign b_s[303308:301800] = s_w_200;
assign b_c[304817:303309] = c_w_201;assign b_s[304817:303309] = s_w_201;
assign b_c[306326:304818] = c_w_202;assign b_s[306326:304818] = s_w_202;
assign b_c[307835:306327] = c_w_203;assign b_s[307835:306327] = s_w_203;
assign b_c[309344:307836] = c_w_204;assign b_s[309344:307836] = s_w_204;
assign b_c[310853:309345] = c_w_205;assign b_s[310853:309345] = s_w_205;
assign b_c[312362:310854] = c_w_206;assign b_s[312362:310854] = s_w_206;
assign b_c[313871:312363] = c_w_207;assign b_s[313871:312363] = s_w_207;
assign b_c[315380:313872] = c_w_208;assign b_s[315380:313872] = s_w_208;
assign b_c[316889:315381] = c_w_209;assign b_s[316889:315381] = s_w_209;
assign b_c[318398:316890] = c_w_210;assign b_s[318398:316890] = s_w_210;
assign b_c[319907:318399] = c_w_211;assign b_s[319907:318399] = s_w_211;
assign b_c[321416:319908] = c_w_212;assign b_s[321416:319908] = s_w_212;
assign b_c[322925:321417] = c_w_213;assign b_s[322925:321417] = s_w_213;
assign b_c[324434:322926] = c_w_214;assign b_s[324434:322926] = s_w_214;
assign b_c[325943:324435] = c_w_215;assign b_s[325943:324435] = s_w_215;
assign b_c[327452:325944] = c_w_216;assign b_s[327452:325944] = s_w_216;
assign b_c[328961:327453] = c_w_217;assign b_s[328961:327453] = s_w_217;
assign b_c[330470:328962] = c_w_218;assign b_s[330470:328962] = s_w_218;
assign b_c[331979:330471] = c_w_219;assign b_s[331979:330471] = s_w_219;
assign b_c[333488:331980] = c_w_220;assign b_s[333488:331980] = s_w_220;
assign b_c[334997:333489] = c_w_221;assign b_s[334997:333489] = s_w_221;
assign b_c[336506:334998] = c_w_222;assign b_s[336506:334998] = s_w_222;
assign b_c[338015:336507] = c_w_223;assign b_s[338015:336507] = s_w_223;
assign b_c[339524:338016] = c_w_224;assign b_s[339524:338016] = s_w_224;
assign b_c[341033:339525] = c_w_225;assign b_s[341033:339525] = s_w_225;
assign b_c[342542:341034] = c_w_226;assign b_s[342542:341034] = s_w_226;
assign b_c[344051:342543] = c_w_227;assign b_s[344051:342543] = s_w_227;
assign b_c[345560:344052] = c_w_228;assign b_s[345560:344052] = s_w_228;
assign b_c[347069:345561] = c_w_229;assign b_s[347069:345561] = s_w_229;
assign b_c[348578:347070] = c_w_230;assign b_s[348578:347070] = s_w_230;
assign b_c[350087:348579] = c_w_231;assign b_s[350087:348579] = s_w_231;
assign b_c[351596:350088] = c_w_232;assign b_s[351596:350088] = s_w_232;
assign b_c[353105:351597] = c_w_233;assign b_s[353105:351597] = s_w_233;
assign b_c[354614:353106] = c_w_234;assign b_s[354614:353106] = s_w_234;
assign b_c[356123:354615] = c_w_235;assign b_s[356123:354615] = s_w_235;
assign b_c[357632:356124] = c_w_236;assign b_s[357632:356124] = s_w_236;
assign b_c[359141:357633] = c_w_237;assign b_s[359141:357633] = s_w_237;
assign b_c[360650:359142] = c_w_238;assign b_s[360650:359142] = s_w_238;
assign b_c[362159:360651] = c_w_239;assign b_s[362159:360651] = s_w_239;
assign b_c[363668:362160] = c_w_240;assign b_s[363668:362160] = s_w_240;
assign b_c[365177:363669] = c_w_241;assign b_s[365177:363669] = s_w_241;
assign b_c[366686:365178] = c_w_242;assign b_s[366686:365178] = s_w_242;
assign b_c[368195:366687] = c_w_243;assign b_s[368195:366687] = s_w_243;
assign b_c[369704:368196] = c_w_244;assign b_s[369704:368196] = s_w_244;
assign b_c[371213:369705] = c_w_245;assign b_s[371213:369705] = s_w_245;
assign b_c[372722:371214] = c_w_246;assign b_s[372722:371214] = s_w_246;
assign b_c[374231:372723] = c_w_247;assign b_s[374231:372723] = s_w_247;
assign b_c[375740:374232] = c_w_248;assign b_s[375740:374232] = s_w_248;
assign b_c[377249:375741] = c_w_249;assign b_s[377249:375741] = s_w_249;
assign b_c[378758:377250] = c_w_250;assign b_s[378758:377250] = s_w_250;
assign b_c[380267:378759] = c_w_251;assign b_s[380267:378759] = s_w_251;
assign b_c[381776:380268] = c_w_252;assign b_s[381776:380268] = s_w_252;
assign b_c[383285:381777] = c_w_253;assign b_s[383285:381777] = s_w_253;
assign b_c[384794:383286] = c_w_254;assign b_s[384794:383286] = s_w_254;
assign b_c[386303:384795] = c_w_255;assign b_s[386303:384795] = s_w_255;
assign b_c[387812:386304] = c_w_256;assign b_s[387812:386304] = s_w_256;
assign b_c[389321:387813] = c_w_257;assign b_s[389321:387813] = s_w_257;
assign b_c[390830:389322] = c_w_258;assign b_s[390830:389322] = s_w_258;
assign b_c[392339:390831] = c_w_259;assign b_s[392339:390831] = s_w_259;
assign b_c[393848:392340] = c_w_260;assign b_s[393848:392340] = s_w_260;
assign b_c[395357:393849] = c_w_261;assign b_s[395357:393849] = s_w_261;
assign b_c[396866:395358] = c_w_262;assign b_s[396866:395358] = s_w_262;
assign b_c[398375:396867] = c_w_263;assign b_s[398375:396867] = s_w_263;
assign b_c[399884:398376] = c_w_264;assign b_s[399884:398376] = s_w_264;
assign b_c[401393:399885] = c_w_265;assign b_s[401393:399885] = s_w_265;
assign b_c[402902:401394] = c_w_266;assign b_s[402902:401394] = s_w_266;
assign b_c[404411:402903] = c_w_267;assign b_s[404411:402903] = s_w_267;
assign b_c[405920:404412] = c_w_268;assign b_s[405920:404412] = s_w_268;
assign b_c[407429:405921] = c_w_269;assign b_s[407429:405921] = s_w_269;
assign b_c[408938:407430] = c_w_270;assign b_s[408938:407430] = s_w_270;
assign b_c[410447:408939] = c_w_271;assign b_s[410447:408939] = s_w_271;
assign b_c[411956:410448] = c_w_272;assign b_s[411956:410448] = s_w_272;
assign b_c[413465:411957] = c_w_273;assign b_s[413465:411957] = s_w_273;
assign b_c[414974:413466] = c_w_274;assign b_s[414974:413466] = s_w_274;
assign b_c[416483:414975] = c_w_275;assign b_s[416483:414975] = s_w_275;
assign b_c[417992:416484] = c_w_276;assign b_s[417992:416484] = s_w_276;
assign b_c[419501:417993] = c_w_277;assign b_s[419501:417993] = s_w_277;
assign b_c[421010:419502] = c_w_278;assign b_s[421010:419502] = s_w_278;
assign b_c[422519:421011] = c_w_279;assign b_s[422519:421011] = s_w_279;
assign b_c[424028:422520] = c_w_280;assign b_s[424028:422520] = s_w_280;
assign b_c[425537:424029] = c_w_281;assign b_s[425537:424029] = s_w_281;
assign b_c[427046:425538] = c_w_282;assign b_s[427046:425538] = s_w_282;
assign b_c[428555:427047] = c_w_283;assign b_s[428555:427047] = s_w_283;
assign b_c[430064:428556] = c_w_284;assign b_s[430064:428556] = s_w_284;
assign b_c[431573:430065] = c_w_285;assign b_s[431573:430065] = s_w_285;
assign b_c[433082:431574] = c_w_286;assign b_s[433082:431574] = s_w_286;
assign b_c[434591:433083] = c_w_287;assign b_s[434591:433083] = s_w_287;
assign b_c[436100:434592] = c_w_288;assign b_s[436100:434592] = s_w_288;
assign b_c[437609:436101] = c_w_289;assign b_s[437609:436101] = s_w_289;
assign b_c[439118:437610] = c_w_290;assign b_s[439118:437610] = s_w_290;
assign b_c[440627:439119] = c_w_291;assign b_s[440627:439119] = s_w_291;
assign b_c[442136:440628] = c_w_292;assign b_s[442136:440628] = s_w_292;
assign b_c[443645:442137] = c_w_293;assign b_s[443645:442137] = s_w_293;
assign b_c[445154:443646] = c_w_294;assign b_s[445154:443646] = s_w_294;
assign b_c[446663:445155] = c_w_295;assign b_s[446663:445155] = s_w_295;
assign b_c[448172:446664] = c_w_296;assign b_s[448172:446664] = s_w_296;
assign b_c[449681:448173] = c_w_297;assign b_s[449681:448173] = s_w_297;
assign b_c[451190:449682] = c_w_298;assign b_s[451190:449682] = s_w_298;
assign b_c[452699:451191] = c_w_299;assign b_s[452699:451191] = s_w_299;
assign b_c[454208:452700] = c_w_300;assign b_s[454208:452700] = s_w_300;
assign b_c[455717:454209] = c_w_301;assign b_s[455717:454209] = s_w_301;
assign b_c[457226:455718] = c_w_302;assign b_s[457226:455718] = s_w_302;
assign b_c[458735:457227] = c_w_303;assign b_s[458735:457227] = s_w_303;
assign b_c[460244:458736] = c_w_304;assign b_s[460244:458736] = s_w_304;
assign b_c[461753:460245] = c_w_305;assign b_s[461753:460245] = s_w_305;
assign b_c[463262:461754] = c_w_306;assign b_s[463262:461754] = s_w_306;
assign b_c[464771:463263] = c_w_307;assign b_s[464771:463263] = s_w_307;
assign b_c[466280:464772] = c_w_308;assign b_s[466280:464772] = s_w_308;
assign b_c[467789:466281] = c_w_309;assign b_s[467789:466281] = s_w_309;
assign b_c[469298:467790] = c_w_310;assign b_s[469298:467790] = s_w_310;
assign b_c[470807:469299] = c_w_311;assign b_s[470807:469299] = s_w_311;
assign b_c[472316:470808] = c_w_312;assign b_s[472316:470808] = s_w_312;
assign b_c[473825:472317] = c_w_313;assign b_s[473825:472317] = s_w_313;
assign b_c[475334:473826] = c_w_314;assign b_s[475334:473826] = s_w_314;
assign b_c[476843:475335] = c_w_315;assign b_s[476843:475335] = s_w_315;
assign b_c[478352:476844] = c_w_316;assign b_s[478352:476844] = s_w_316;
assign b_c[479861:478353] = c_w_317;assign b_s[479861:478353] = s_w_317;
assign b_c[481370:479862] = c_w_318;assign b_s[481370:479862] = s_w_318;
assign b_c[482879:481371] = c_w_319;assign b_s[482879:481371] = s_w_319;
assign b_c[484388:482880] = c_w_320;assign b_s[484388:482880] = s_w_320;
assign b_c[485897:484389] = c_w_321;assign b_s[485897:484389] = s_w_321;
assign b_c[487406:485898] = c_w_322;assign b_s[487406:485898] = s_w_322;
assign b_c[488915:487407] = c_w_323;assign b_s[488915:487407] = s_w_323;
assign b_c[490424:488916] = c_w_324;assign b_s[490424:488916] = s_w_324;
assign b_c[491933:490425] = c_w_325;assign b_s[491933:490425] = s_w_325;
assign b_c[493442:491934] = c_w_326;assign b_s[493442:491934] = s_w_326;
assign b_c[494951:493443] = c_w_327;assign b_s[494951:493443] = s_w_327;
assign b_c[496460:494952] = c_w_328;assign b_s[496460:494952] = s_w_328;
assign b_c[497969:496461] = c_w_329;assign b_s[497969:496461] = s_w_329;
assign b_c[499478:497970] = c_w_330;assign b_s[499478:497970] = s_w_330;
assign b_c[500987:499479] = c_w_331;assign b_s[500987:499479] = s_w_331;
assign b_c[502496:500988] = c_w_332;assign b_s[502496:500988] = s_w_332;
assign b_c[504005:502497] = c_w_333;assign b_s[504005:502497] = s_w_333;
assign b_c[505514:504006] = c_w_334;assign b_s[505514:504006] = s_w_334;
assign b_c[507023:505515] = c_w_335;assign b_s[507023:505515] = s_w_335;
assign b_c[508532:507024] = c_w_336;assign b_s[508532:507024] = s_w_336;
assign b_c[510041:508533] = c_w_337;assign b_s[510041:508533] = s_w_337;
assign b_c[511550:510042] = c_w_338;assign b_s[511550:510042] = s_w_338;
assign b_c[513059:511551] = c_w_339;assign b_s[513059:511551] = s_w_339;
assign b_c[514568:513060] = c_w_340;assign b_s[514568:513060] = s_w_340;
assign b_c[516077:514569] = c_w_341;assign b_s[516077:514569] = s_w_341;
assign b_c[517586:516078] = c_w_342;assign b_s[517586:516078] = s_w_342;
assign b_c[519095:517587] = c_w_343;assign b_s[519095:517587] = s_w_343;
assign b_c[520604:519096] = c_w_344;assign b_s[520604:519096] = s_w_344;
assign b_c[522113:520605] = c_w_345;assign b_s[522113:520605] = s_w_345;
assign b_c[523622:522114] = c_w_346;assign b_s[523622:522114] = s_w_346;
assign b_c[525131:523623] = c_w_347;assign b_s[525131:523623] = s_w_347;
assign b_c[526640:525132] = c_w_348;assign b_s[526640:525132] = s_w_348;
assign b_c[528149:526641] = c_w_349;assign b_s[528149:526641] = s_w_349;
assign b_c[529658:528150] = c_w_350;assign b_s[529658:528150] = s_w_350;
assign b_c[531167:529659] = c_w_351;assign b_s[531167:529659] = s_w_351;
assign b_c[532676:531168] = c_w_352;assign b_s[532676:531168] = s_w_352;
assign b_c[534185:532677] = c_w_353;assign b_s[534185:532677] = s_w_353;
assign b_c[535694:534186] = c_w_354;assign b_s[535694:534186] = s_w_354;
assign b_c[537203:535695] = c_w_355;assign b_s[537203:535695] = s_w_355;
assign b_c[538712:537204] = c_w_356;assign b_s[538712:537204] = s_w_356;
assign b_c[540221:538713] = c_w_357;assign b_s[540221:538713] = s_w_357;
assign b_c[541730:540222] = c_w_358;assign b_s[541730:540222] = s_w_358;
assign b_c[543239:541731] = c_w_359;assign b_s[543239:541731] = s_w_359;
assign b_c[544748:543240] = c_w_360;assign b_s[544748:543240] = s_w_360;
assign b_c[546257:544749] = c_w_361;assign b_s[546257:544749] = s_w_361;
assign b_c[547766:546258] = c_w_362;assign b_s[547766:546258] = s_w_362;
assign b_c[549275:547767] = c_w_363;assign b_s[549275:547767] = s_w_363;
assign b_c[550784:549276] = c_w_364;assign b_s[550784:549276] = s_w_364;
assign b_c[552293:550785] = c_w_365;assign b_s[552293:550785] = s_w_365;
assign b_c[553802:552294] = c_w_366;assign b_s[553802:552294] = s_w_366;
assign b_c[555311:553803] = c_w_367;assign b_s[555311:553803] = s_w_367;
assign b_c[556820:555312] = c_w_368;assign b_s[556820:555312] = s_w_368;
assign b_c[558329:556821] = c_w_369;assign b_s[558329:556821] = s_w_369;
assign b_c[559838:558330] = c_w_370;assign b_s[559838:558330] = s_w_370;
assign b_c[561347:559839] = c_w_371;assign b_s[561347:559839] = s_w_371;
assign b_c[562856:561348] = c_w_372;assign b_s[562856:561348] = s_w_372;
assign b_c[564365:562857] = c_w_373;assign b_s[564365:562857] = s_w_373;
assign b_c[565874:564366] = c_w_374;assign b_s[565874:564366] = s_w_374;
assign b_c[567383:565875] = c_w_375;assign b_s[567383:565875] = s_w_375;
assign b_c[568892:567384] = c_w_376;assign b_s[568892:567384] = s_w_376;
assign b_c[570401:568893] = c_w_377;assign b_s[570401:568893] = s_w_377;
assign b_c[571910:570402] = c_w_378;assign b_s[571910:570402] = s_w_378;
assign b_c[573419:571911] = c_w_379;assign b_s[573419:571911] = s_w_379;
assign b_c[574928:573420] = c_w_380;assign b_s[574928:573420] = s_w_380;
assign b_c[576437:574929] = c_w_381;assign b_s[576437:574929] = s_w_381;
assign b_c[577946:576438] = c_w_382;assign b_s[577946:576438] = s_w_382;
assign b_c[579455:577947] = c_w_383;assign b_s[579455:577947] = s_w_383;
assign b_c[580964:579456] = c_w_384;assign b_s[580964:579456] = s_w_384;
assign b_c[582473:580965] = c_w_385;assign b_s[582473:580965] = s_w_385;
assign b_c[583982:582474] = c_w_386;assign b_s[583982:582474] = s_w_386;
assign b_c[585491:583983] = c_w_387;assign b_s[585491:583983] = s_w_387;
assign b_c[587000:585492] = c_w_388;assign b_s[587000:585492] = s_w_388;
assign b_c[588509:587001] = c_w_389;assign b_s[588509:587001] = s_w_389;
assign b_c[590018:588510] = c_w_390;assign b_s[590018:588510] = s_w_390;
assign b_c[591527:590019] = c_w_391;assign b_s[591527:590019] = s_w_391;
assign b_c[593036:591528] = c_w_392;assign b_s[593036:591528] = s_w_392;
assign b_c[594545:593037] = c_w_393;assign b_s[594545:593037] = s_w_393;
assign b_c[596054:594546] = c_w_394;assign b_s[596054:594546] = s_w_394;
assign b_c[597563:596055] = c_w_395;assign b_s[597563:596055] = s_w_395;
assign b_c[599072:597564] = c_w_396;assign b_s[599072:597564] = s_w_396;
assign b_c[600581:599073] = c_w_397;assign b_s[600581:599073] = s_w_397;
assign b_c[602090:600582] = c_w_398;assign b_s[602090:600582] = s_w_398;
assign b_c[603599:602091] = c_w_399;assign b_s[603599:602091] = s_w_399;
assign b_c[605108:603600] = c_w_400;assign b_s[605108:603600] = s_w_400;
assign b_c[606617:605109] = c_w_401;assign b_s[606617:605109] = s_w_401;
assign b_c[608126:606618] = c_w_402;assign b_s[608126:606618] = s_w_402;
assign b_c[609635:608127] = c_w_403;assign b_s[609635:608127] = s_w_403;
assign b_c[611144:609636] = c_w_404;assign b_s[611144:609636] = s_w_404;
assign b_c[612653:611145] = c_w_405;assign b_s[612653:611145] = s_w_405;
assign b_c[614162:612654] = c_w_406;assign b_s[614162:612654] = s_w_406;
assign b_c[615671:614163] = c_w_407;assign b_s[615671:614163] = s_w_407;
assign b_c[617180:615672] = c_w_408;assign b_s[617180:615672] = s_w_408;
assign b_c[618689:617181] = c_w_409;assign b_s[618689:617181] = s_w_409;
assign b_c[620198:618690] = c_w_410;assign b_s[620198:618690] = s_w_410;
assign b_c[621707:620199] = c_w_411;assign b_s[621707:620199] = s_w_411;
assign b_c[623216:621708] = c_w_412;assign b_s[623216:621708] = s_w_412;
assign b_c[624725:623217] = c_w_413;assign b_s[624725:623217] = s_w_413;
assign b_c[626234:624726] = c_w_414;assign b_s[626234:624726] = s_w_414;
assign b_c[627743:626235] = c_w_415;assign b_s[627743:626235] = s_w_415;
assign b_c[629252:627744] = c_w_416;assign b_s[629252:627744] = s_w_416;
assign b_c[630761:629253] = c_w_417;assign b_s[630761:629253] = s_w_417;
assign b_c[632270:630762] = c_w_418;assign b_s[632270:630762] = s_w_418;
assign b_c[633779:632271] = c_w_419;assign b_s[633779:632271] = s_w_419;
assign b_c[635288:633780] = c_w_420;assign b_s[635288:633780] = s_w_420;
assign b_c[636797:635289] = c_w_421;assign b_s[636797:635289] = s_w_421;
assign b_c[638306:636798] = c_w_422;assign b_s[638306:636798] = s_w_422;
assign b_c[639815:638307] = c_w_423;assign b_s[639815:638307] = s_w_423;
assign b_c[641324:639816] = c_w_424;assign b_s[641324:639816] = s_w_424;
assign b_c[642833:641325] = c_w_425;assign b_s[642833:641325] = s_w_425;
assign b_c[644342:642834] = c_w_426;assign b_s[644342:642834] = s_w_426;
assign b_c[645851:644343] = c_w_427;assign b_s[645851:644343] = s_w_427;
assign b_c[647360:645852] = c_w_428;assign b_s[647360:645852] = s_w_428;
assign b_c[648869:647361] = c_w_429;assign b_s[648869:647361] = s_w_429;
assign b_c[650378:648870] = c_w_430;assign b_s[650378:648870] = s_w_430;
assign b_c[651887:650379] = c_w_431;assign b_s[651887:650379] = s_w_431;
assign b_c[653396:651888] = c_w_432;assign b_s[653396:651888] = s_w_432;
assign b_c[654905:653397] = c_w_433;assign b_s[654905:653397] = s_w_433;
assign b_c[656414:654906] = c_w_434;assign b_s[656414:654906] = s_w_434;
assign b_c[657923:656415] = c_w_435;assign b_s[657923:656415] = s_w_435;
assign b_c[659432:657924] = c_w_436;assign b_s[659432:657924] = s_w_436;
assign b_c[660941:659433] = c_w_437;assign b_s[660941:659433] = s_w_437;
assign b_c[662450:660942] = c_w_438;assign b_s[662450:660942] = s_w_438;
assign b_c[663959:662451] = c_w_439;assign b_s[663959:662451] = s_w_439;
assign b_c[665468:663960] = c_w_440;assign b_s[665468:663960] = s_w_440;
assign b_c[666977:665469] = c_w_441;assign b_s[666977:665469] = s_w_441;
assign b_c[668486:666978] = c_w_442;assign b_s[668486:666978] = s_w_442;
assign b_c[669995:668487] = c_w_443;assign b_s[669995:668487] = s_w_443;
assign b_c[671504:669996] = c_w_444;assign b_s[671504:669996] = s_w_444;
assign b_c[673013:671505] = c_w_445;assign b_s[673013:671505] = s_w_445;
assign b_c[674522:673014] = c_w_446;assign b_s[674522:673014] = s_w_446;
assign b_c[676031:674523] = c_w_447;assign b_s[676031:674523] = s_w_447;
assign b_c[677540:676032] = c_w_448;assign b_s[677540:676032] = s_w_448;
assign b_c[679049:677541] = c_w_449;assign b_s[679049:677541] = s_w_449;
assign b_c[680558:679050] = c_w_450;assign b_s[680558:679050] = s_w_450;
assign b_c[682067:680559] = c_w_451;assign b_s[682067:680559] = s_w_451;
assign b_c[683576:682068] = c_w_452;assign b_s[683576:682068] = s_w_452;
assign b_c[685085:683577] = c_w_453;assign b_s[685085:683577] = s_w_453;
assign b_c[686594:685086] = c_w_454;assign b_s[686594:685086] = s_w_454;
assign b_c[688103:686595] = c_w_455;assign b_s[688103:686595] = s_w_455;
assign b_c[689612:688104] = c_w_456;assign b_s[689612:688104] = s_w_456;
assign b_c[691121:689613] = c_w_457;assign b_s[691121:689613] = s_w_457;
assign b_c[692630:691122] = c_w_458;assign b_s[692630:691122] = s_w_458;
assign b_c[694139:692631] = c_w_459;assign b_s[694139:692631] = s_w_459;
assign b_c[695648:694140] = c_w_460;assign b_s[695648:694140] = s_w_460;
assign b_c[697157:695649] = c_w_461;assign b_s[697157:695649] = s_w_461;
assign b_c[698666:697158] = c_w_462;assign b_s[698666:697158] = s_w_462;
assign b_c[700175:698667] = c_w_463;assign b_s[700175:698667] = s_w_463;
assign b_c[701684:700176] = c_w_464;assign b_s[701684:700176] = s_w_464;
assign b_c[703193:701685] = c_w_465;assign b_s[703193:701685] = s_w_465;
assign b_c[704702:703194] = c_w_466;assign b_s[704702:703194] = s_w_466;
assign b_c[706211:704703] = c_w_467;assign b_s[706211:704703] = s_w_467;
assign b_c[707720:706212] = c_w_468;assign b_s[707720:706212] = s_w_468;
assign b_c[709229:707721] = c_w_469;assign b_s[709229:707721] = s_w_469;
assign b_c[710738:709230] = c_w_470;assign b_s[710738:709230] = s_w_470;
assign b_c[712247:710739] = c_w_471;assign b_s[712247:710739] = s_w_471;
assign b_c[713756:712248] = c_w_472;assign b_s[713756:712248] = s_w_472;
assign b_c[715265:713757] = c_w_473;assign b_s[715265:713757] = s_w_473;
assign b_c[716774:715266] = c_w_474;assign b_s[716774:715266] = s_w_474;
assign b_c[718283:716775] = c_w_475;assign b_s[718283:716775] = s_w_475;
assign b_c[719792:718284] = c_w_476;assign b_s[719792:718284] = s_w_476;
assign b_c[721301:719793] = c_w_477;assign b_s[721301:719793] = s_w_477;
assign b_c[722810:721302] = c_w_478;assign b_s[722810:721302] = s_w_478;
assign b_c[724319:722811] = c_w_479;assign b_s[724319:722811] = s_w_479;
assign b_c[725828:724320] = c_w_480;assign b_s[725828:724320] = s_w_480;
assign b_c[727337:725829] = c_w_481;assign b_s[727337:725829] = s_w_481;
assign b_c[728846:727338] = c_w_482;assign b_s[728846:727338] = s_w_482;
assign b_c[730355:728847] = c_w_483;assign b_s[730355:728847] = s_w_483;
assign b_c[731864:730356] = c_w_484;assign b_s[731864:730356] = s_w_484;
assign b_c[733373:731865] = c_w_485;assign b_s[733373:731865] = s_w_485;
assign b_c[734882:733374] = c_w_486;assign b_s[734882:733374] = s_w_486;
assign b_c[736391:734883] = c_w_487;assign b_s[736391:734883] = s_w_487;
assign b_c[737900:736392] = c_w_488;assign b_s[737900:736392] = s_w_488;
assign b_c[739409:737901] = c_w_489;assign b_s[739409:737901] = s_w_489;
assign b_c[740918:739410] = c_w_490;assign b_s[740918:739410] = s_w_490;
assign b_c[742427:740919] = c_w_491;assign b_s[742427:740919] = s_w_491;
assign b_c[743936:742428] = c_w_492;assign b_s[743936:742428] = s_w_492;
assign b_c[745445:743937] = c_w_493;assign b_s[745445:743937] = s_w_493;
assign b_c[746954:745446] = c_w_494;assign b_s[746954:745446] = s_w_494;
assign b_c[748463:746955] = c_w_495;assign b_s[748463:746955] = s_w_495;
assign b_c[749972:748464] = c_w_496;assign b_s[749972:748464] = s_w_496;
assign b_c[751481:749973] = c_w_497;assign b_s[751481:749973] = s_w_497;
assign b_c[752990:751482] = c_w_498;assign b_s[752990:751482] = s_w_498;
assign b_c[754499:752991] = c_w_499;assign b_s[754499:752991] = s_w_499;
assign b_c[756008:754500] = c_w_500;assign b_s[756008:754500] = s_w_500;
assign b_c[757517:756009] = c_w_501;assign b_s[757517:756009] = s_w_501;
assign b_c[759026:757518] = c_w_502;assign b_s[759026:757518] = s_w_502;
assign b_c[760535:759027] = c_w_503;assign b_s[760535:759027] = s_w_503;
assign b_c[762044:760536] = c_w_504;assign b_s[762044:760536] = s_w_504;
assign b_c[763553:762045] = c_w_505;assign b_s[763553:762045] = s_w_505;
assign b_c[765062:763554] = c_w_506;assign b_s[765062:763554] = s_w_506;
assign b_c[766571:765063] = c_w_507;assign b_s[766571:765063] = s_w_507;
assign b_c[768080:766572] = c_w_508;assign b_s[768080:766572] = s_w_508;
assign b_c[769589:768081] = c_w_509;assign b_s[769589:768081] = s_w_509;
assign b_c[771098:769590] = c_w_510;assign b_s[771098:769590] = s_w_510;
assign b_c[772607:771099] = c_w_511;assign b_s[772607:771099] = s_w_511;
assign b_c[774116:772608] = c_w_512;assign b_s[774116:772608] = s_w_512;
assign b_c[775625:774117] = c_w_513;assign b_s[775625:774117] = s_w_513;
assign b_c[777134:775626] = c_w_514;assign b_s[777134:775626] = s_w_514;
assign b_c[778643:777135] = c_w_515;assign b_s[778643:777135] = s_w_515;
assign b_c[780152:778644] = c_w_516;assign b_s[780152:778644] = s_w_516;
assign b_c[781661:780153] = c_w_517;assign b_s[781661:780153] = s_w_517;
assign b_c[783170:781662] = c_w_518;assign b_s[783170:781662] = s_w_518;
assign b_c[784679:783171] = c_w_519;assign b_s[784679:783171] = s_w_519;
assign b_c[786188:784680] = c_w_520;assign b_s[786188:784680] = s_w_520;
assign b_c[787697:786189] = c_w_521;assign b_s[787697:786189] = s_w_521;
assign b_c[789206:787698] = c_w_522;assign b_s[789206:787698] = s_w_522;
assign b_c[790715:789207] = c_w_523;assign b_s[790715:789207] = s_w_523;
assign b_c[792224:790716] = c_w_524;assign b_s[792224:790716] = s_w_524;
assign b_c[793733:792225] = c_w_525;assign b_s[793733:792225] = s_w_525;
assign b_c[795242:793734] = c_w_526;assign b_s[795242:793734] = s_w_526;
assign b_c[796751:795243] = c_w_527;assign b_s[796751:795243] = s_w_527;
assign b_c[798260:796752] = c_w_528;assign b_s[798260:796752] = s_w_528;
assign b_c[799769:798261] = c_w_529;assign b_s[799769:798261] = s_w_529;
assign b_c[801278:799770] = c_w_530;assign b_s[801278:799770] = s_w_530;
assign b_c[802787:801279] = c_w_531;assign b_s[802787:801279] = s_w_531;
assign b_c[804296:802788] = c_w_532;assign b_s[804296:802788] = s_w_532;
assign b_c[805805:804297] = c_w_533;assign b_s[805805:804297] = s_w_533;
assign b_c[807314:805806] = c_w_534;assign b_s[807314:805806] = s_w_534;
assign b_c[808823:807315] = c_w_535;assign b_s[808823:807315] = s_w_535;
assign b_c[810332:808824] = c_w_536;assign b_s[810332:808824] = s_w_536;
assign b_c[811841:810333] = c_w_537;assign b_s[811841:810333] = s_w_537;
assign b_c[813350:811842] = c_w_538;assign b_s[813350:811842] = s_w_538;
assign b_c[814859:813351] = c_w_539;assign b_s[814859:813351] = s_w_539;
assign b_c[816368:814860] = c_w_540;assign b_s[816368:814860] = s_w_540;
assign b_c[817877:816369] = c_w_541;assign b_s[817877:816369] = s_w_541;
assign b_c[819386:817878] = c_w_542;assign b_s[819386:817878] = s_w_542;
assign b_c[820895:819387] = c_w_543;assign b_s[820895:819387] = s_w_543;
assign b_c[822404:820896] = c_w_544;assign b_s[822404:820896] = s_w_544;
assign b_c[823913:822405] = c_w_545;assign b_s[823913:822405] = s_w_545;
assign b_c[825422:823914] = c_w_546;assign b_s[825422:823914] = s_w_546;
assign b_c[826931:825423] = c_w_547;assign b_s[826931:825423] = s_w_547;
assign b_c[828440:826932] = c_w_548;assign b_s[828440:826932] = s_w_548;
assign b_c[829949:828441] = c_w_549;assign b_s[829949:828441] = s_w_549;
assign b_c[831458:829950] = c_w_550;assign b_s[831458:829950] = s_w_550;
assign b_c[832967:831459] = c_w_551;assign b_s[832967:831459] = s_w_551;
assign b_c[834476:832968] = c_w_552;assign b_s[834476:832968] = s_w_552;
assign b_c[835985:834477] = c_w_553;assign b_s[835985:834477] = s_w_553;
assign b_c[837494:835986] = c_w_554;assign b_s[837494:835986] = s_w_554;
assign b_c[839003:837495] = c_w_555;assign b_s[839003:837495] = s_w_555;
assign b_c[840512:839004] = c_w_556;assign b_s[840512:839004] = s_w_556;
assign b_c[842021:840513] = c_w_557;assign b_s[842021:840513] = s_w_557;
assign b_c[843530:842022] = c_w_558;assign b_s[843530:842022] = s_w_558;
assign b_c[845039:843531] = c_w_559;assign b_s[845039:843531] = s_w_559;
assign b_c[846548:845040] = c_w_560;assign b_s[846548:845040] = s_w_560;
assign b_c[848057:846549] = c_w_561;assign b_s[848057:846549] = s_w_561;
assign b_c[849566:848058] = c_w_562;assign b_s[849566:848058] = s_w_562;
assign b_c[851075:849567] = c_w_563;assign b_s[851075:849567] = s_w_563;
assign b_c[852584:851076] = c_w_564;assign b_s[852584:851076] = s_w_564;
assign b_c[854093:852585] = c_w_565;assign b_s[854093:852585] = s_w_565;
assign b_c[855602:854094] = c_w_566;assign b_s[855602:854094] = s_w_566;
assign b_c[857111:855603] = c_w_567;assign b_s[857111:855603] = s_w_567;
assign b_c[858620:857112] = c_w_568;assign b_s[858620:857112] = s_w_568;
assign b_c[860129:858621] = c_w_569;assign b_s[860129:858621] = s_w_569;
assign b_c[861638:860130] = c_w_570;assign b_s[861638:860130] = s_w_570;
assign b_c[863147:861639] = c_w_571;assign b_s[863147:861639] = s_w_571;
assign b_c[864656:863148] = c_w_572;assign b_s[864656:863148] = s_w_572;
assign b_c[866165:864657] = c_w_573;assign b_s[866165:864657] = s_w_573;
assign b_c[867674:866166] = c_w_574;assign b_s[867674:866166] = s_w_574;
assign b_c[869183:867675] = c_w_575;assign b_s[869183:867675] = s_w_575;
assign b_c[870692:869184] = c_w_576;assign b_s[870692:869184] = s_w_576;
assign b_c[872201:870693] = c_w_577;assign b_s[872201:870693] = s_w_577;
assign b_c[873710:872202] = c_w_578;assign b_s[873710:872202] = s_w_578;
assign b_c[875219:873711] = c_w_579;assign b_s[875219:873711] = s_w_579;
assign b_c[876728:875220] = c_w_580;assign b_s[876728:875220] = s_w_580;
assign b_c[878237:876729] = c_w_581;assign b_s[878237:876729] = s_w_581;
assign b_c[879746:878238] = c_w_582;assign b_s[879746:878238] = s_w_582;
assign b_c[881255:879747] = c_w_583;assign b_s[881255:879747] = s_w_583;
assign b_c[882764:881256] = c_w_584;assign b_s[882764:881256] = s_w_584;
assign b_c[884273:882765] = c_w_585;assign b_s[884273:882765] = s_w_585;
assign b_c[885782:884274] = c_w_586;assign b_s[885782:884274] = s_w_586;
assign b_c[887291:885783] = c_w_587;assign b_s[887291:885783] = s_w_587;
assign b_c[888800:887292] = c_w_588;assign b_s[888800:887292] = s_w_588;
assign b_c[890309:888801] = c_w_589;assign b_s[890309:888801] = s_w_589;
assign b_c[891818:890310] = c_w_590;assign b_s[891818:890310] = s_w_590;
assign b_c[893327:891819] = c_w_591;assign b_s[893327:891819] = s_w_591;
assign b_c[894836:893328] = c_w_592;assign b_s[894836:893328] = s_w_592;
assign b_c[896345:894837] = c_w_593;assign b_s[896345:894837] = s_w_593;
assign b_c[897854:896346] = c_w_594;assign b_s[897854:896346] = s_w_594;
assign b_c[899363:897855] = c_w_595;assign b_s[899363:897855] = s_w_595;
assign b_c[900872:899364] = c_w_596;assign b_s[900872:899364] = s_w_596;
assign b_c[902381:900873] = c_w_597;assign b_s[902381:900873] = s_w_597;
assign b_c[903890:902382] = c_w_598;assign b_s[903890:902382] = s_w_598;
assign b_c[905399:903891] = c_w_599;assign b_s[905399:903891] = s_w_599;
assign b_c[906908:905400] = c_w_600;assign b_s[906908:905400] = s_w_600;
assign b_c[908417:906909] = c_w_601;assign b_s[908417:906909] = s_w_601;
assign b_c[909926:908418] = c_w_602;assign b_s[909926:908418] = s_w_602;
assign b_c[911435:909927] = c_w_603;assign b_s[911435:909927] = s_w_603;
assign b_c[912944:911436] = c_w_604;assign b_s[912944:911436] = s_w_604;
assign b_c[914453:912945] = c_w_605;assign b_s[914453:912945] = s_w_605;
assign b_c[915962:914454] = c_w_606;assign b_s[915962:914454] = s_w_606;
assign b_c[917471:915963] = c_w_607;assign b_s[917471:915963] = s_w_607;
assign b_c[918980:917472] = c_w_608;assign b_s[918980:917472] = s_w_608;
assign b_c[920489:918981] = c_w_609;assign b_s[920489:918981] = s_w_609;
assign b_c[921998:920490] = c_w_610;assign b_s[921998:920490] = s_w_610;
assign b_c[923507:921999] = c_w_611;assign b_s[923507:921999] = s_w_611;
assign b_c[925016:923508] = c_w_612;assign b_s[925016:923508] = s_w_612;
assign b_c[926525:925017] = c_w_613;assign b_s[926525:925017] = s_w_613;
assign b_c[928034:926526] = c_w_614;assign b_s[928034:926526] = s_w_614;
assign b_c[929543:928035] = c_w_615;assign b_s[929543:928035] = s_w_615;
assign b_c[931052:929544] = c_w_616;assign b_s[931052:929544] = s_w_616;
assign b_c[932561:931053] = c_w_617;assign b_s[932561:931053] = s_w_617;
assign b_c[934070:932562] = c_w_618;assign b_s[934070:932562] = s_w_618;
assign b_c[935579:934071] = c_w_619;assign b_s[935579:934071] = s_w_619;
assign b_c[937088:935580] = c_w_620;assign b_s[937088:935580] = s_w_620;
assign b_c[938597:937089] = c_w_621;assign b_s[938597:937089] = s_w_621;
assign b_c[940106:938598] = c_w_622;assign b_s[940106:938598] = s_w_622;
assign b_c[941615:940107] = c_w_623;assign b_s[941615:940107] = s_w_623;
assign b_c[943124:941616] = c_w_624;assign b_s[943124:941616] = s_w_624;
assign b_c[944633:943125] = c_w_625;assign b_s[944633:943125] = s_w_625;
assign b_c[946142:944634] = c_w_626;assign b_s[946142:944634] = s_w_626;
assign b_c[947651:946143] = c_w_627;assign b_s[947651:946143] = s_w_627;
assign b_c[949160:947652] = c_w_628;assign b_s[949160:947652] = s_w_628;
assign b_c[950669:949161] = c_w_629;assign b_s[950669:949161] = s_w_629;
assign b_c[952178:950670] = c_w_630;assign b_s[952178:950670] = s_w_630;
assign b_c[953687:952179] = c_w_631;assign b_s[953687:952179] = s_w_631;
assign b_c[955196:953688] = c_w_632;assign b_s[955196:953688] = s_w_632;
assign b_c[956705:955197] = c_w_633;assign b_s[956705:955197] = s_w_633;
assign b_c[958214:956706] = c_w_634;assign b_s[958214:956706] = s_w_634;
assign b_c[959723:958215] = c_w_635;assign b_s[959723:958215] = s_w_635;
assign b_c[961232:959724] = c_w_636;assign b_s[961232:959724] = s_w_636;
assign b_c[962741:961233] = c_w_637;assign b_s[962741:961233] = s_w_637;
assign b_c[964250:962742] = c_w_638;assign b_s[964250:962742] = s_w_638;
assign b_c[965759:964251] = c_w_639;assign b_s[965759:964251] = s_w_639;
assign b_c[967268:965760] = c_w_640;assign b_s[967268:965760] = s_w_640;
assign b_c[968777:967269] = c_w_641;assign b_s[968777:967269] = s_w_641;
assign b_c[970286:968778] = c_w_642;assign b_s[970286:968778] = s_w_642;
assign b_c[971795:970287] = c_w_643;assign b_s[971795:970287] = s_w_643;
assign b_c[973304:971796] = c_w_644;assign b_s[973304:971796] = s_w_644;
assign b_c[974813:973305] = c_w_645;assign b_s[974813:973305] = s_w_645;
assign b_c[976322:974814] = c_w_646;assign b_s[976322:974814] = s_w_646;
assign b_c[977831:976323] = c_w_647;assign b_s[977831:976323] = s_w_647;
assign b_c[979340:977832] = c_w_648;assign b_s[979340:977832] = s_w_648;
assign b_c[980849:979341] = c_w_649;assign b_s[980849:979341] = s_w_649;
assign b_c[982358:980850] = c_w_650;assign b_s[982358:980850] = s_w_650;
assign b_c[983867:982359] = c_w_651;assign b_s[983867:982359] = s_w_651;
assign b_c[985376:983868] = c_w_652;assign b_s[985376:983868] = s_w_652;
assign b_c[986885:985377] = c_w_653;assign b_s[986885:985377] = s_w_653;
assign b_c[988394:986886] = c_w_654;assign b_s[988394:986886] = s_w_654;
assign b_c[989903:988395] = c_w_655;assign b_s[989903:988395] = s_w_655;
assign b_c[991412:989904] = c_w_656;assign b_s[991412:989904] = s_w_656;
assign b_c[992921:991413] = c_w_657;assign b_s[992921:991413] = s_w_657;
assign b_c[994430:992922] = c_w_658;assign b_s[994430:992922] = s_w_658;
assign b_c[995939:994431] = c_w_659;assign b_s[995939:994431] = s_w_659;
assign b_c[997448:995940] = c_w_660;assign b_s[997448:995940] = s_w_660;
assign b_c[998957:997449] = c_w_661;assign b_s[998957:997449] = s_w_661;
assign b_c[1000466:998958] = c_w_662;assign b_s[1000466:998958] = s_w_662;
assign b_c[1001975:1000467] = c_w_663;assign b_s[1001975:1000467] = s_w_663;
assign b_c[1003484:1001976] = c_w_664;assign b_s[1003484:1001976] = s_w_664;
assign b_c[1004993:1003485] = c_w_665;assign b_s[1004993:1003485] = s_w_665;
assign b_c[1006502:1004994] = c_w_666;assign b_s[1006502:1004994] = s_w_666;
assign b_c[1008011:1006503] = c_w_667;assign b_s[1008011:1006503] = s_w_667;
assign b_c[1009520:1008012] = c_w_668;assign b_s[1009520:1008012] = s_w_668;
assign b_c[1011029:1009521] = c_w_669;assign b_s[1011029:1009521] = s_w_669;
assign b_c[1012538:1011030] = c_w_670;assign b_s[1012538:1011030] = s_w_670;
assign b_c[1014047:1012539] = c_w_671;assign b_s[1014047:1012539] = s_w_671;
assign b_c[1015556:1014048] = c_w_672;assign b_s[1015556:1014048] = s_w_672;
assign b_c[1017065:1015557] = c_w_673;assign b_s[1017065:1015557] = s_w_673;
assign b_c[1018574:1017066] = c_w_674;assign b_s[1018574:1017066] = s_w_674;
assign b_c[1020083:1018575] = c_w_675;assign b_s[1020083:1018575] = s_w_675;
assign b_c[1021592:1020084] = c_w_676;assign b_s[1021592:1020084] = s_w_676;
assign b_c[1023101:1021593] = c_w_677;assign b_s[1023101:1021593] = s_w_677;
assign b_c[1024610:1023102] = c_w_678;assign b_s[1024610:1023102] = s_w_678;
assign b_c[1026119:1024611] = c_w_679;assign b_s[1026119:1024611] = s_w_679;
assign b_c[1027628:1026120] = c_w_680;assign b_s[1027628:1026120] = s_w_680;
assign b_c[1029137:1027629] = c_w_681;assign b_s[1029137:1027629] = s_w_681;
assign b_c[1030646:1029138] = c_w_682;assign b_s[1030646:1029138] = s_w_682;
assign b_c[1032155:1030647] = c_w_683;assign b_s[1032155:1030647] = s_w_683;
assign b_c[1033664:1032156] = c_w_684;assign b_s[1033664:1032156] = s_w_684;
assign b_c[1035173:1033665] = c_w_685;assign b_s[1035173:1033665] = s_w_685;
assign b_c[1036682:1035174] = c_w_686;assign b_s[1036682:1035174] = s_w_686;
assign b_c[1038191:1036683] = c_w_687;assign b_s[1038191:1036683] = s_w_687;
assign b_c[1039700:1038192] = c_w_688;assign b_s[1039700:1038192] = s_w_688;
assign b_c[1041209:1039701] = c_w_689;assign b_s[1041209:1039701] = s_w_689;
assign b_c[1042718:1041210] = c_w_690;assign b_s[1042718:1041210] = s_w_690;
assign b_c[1044227:1042719] = c_w_691;assign b_s[1044227:1042719] = s_w_691;
assign b_c[1045736:1044228] = c_w_692;assign b_s[1045736:1044228] = s_w_692;
assign b_c[1047245:1045737] = c_w_693;assign b_s[1047245:1045737] = s_w_693;
assign b_c[1048754:1047246] = c_w_694;assign b_s[1048754:1047246] = s_w_694;
assign b_c[1050263:1048755] = c_w_695;assign b_s[1050263:1048755] = s_w_695;
assign b_c[1051772:1050264] = c_w_696;assign b_s[1051772:1050264] = s_w_696;
assign b_c[1053281:1051773] = c_w_697;assign b_s[1053281:1051773] = s_w_697;
assign b_c[1054790:1053282] = c_w_698;assign b_s[1054790:1053282] = s_w_698;
assign b_c[1056299:1054791] = c_w_699;assign b_s[1056299:1054791] = s_w_699;
assign b_c[1057808:1056300] = c_w_700;assign b_s[1057808:1056300] = s_w_700;
assign b_c[1059317:1057809] = c_w_701;assign b_s[1059317:1057809] = s_w_701;
assign b_c[1060826:1059318] = c_w_702;assign b_s[1060826:1059318] = s_w_702;
assign b_c[1062335:1060827] = c_w_703;assign b_s[1062335:1060827] = s_w_703;
assign b_c[1063844:1062336] = c_w_704;assign b_s[1063844:1062336] = s_w_704;
assign b_c[1065353:1063845] = c_w_705;assign b_s[1065353:1063845] = s_w_705;
assign b_c[1066862:1065354] = c_w_706;assign b_s[1066862:1065354] = s_w_706;
assign b_c[1068371:1066863] = c_w_707;assign b_s[1068371:1066863] = s_w_707;
assign b_c[1069880:1068372] = c_w_708;assign b_s[1069880:1068372] = s_w_708;
assign b_c[1071389:1069881] = c_w_709;assign b_s[1071389:1069881] = s_w_709;
assign b_c[1072898:1071390] = c_w_710;assign b_s[1072898:1071390] = s_w_710;
assign b_c[1074407:1072899] = c_w_711;assign b_s[1074407:1072899] = s_w_711;
assign b_c[1075916:1074408] = c_w_712;assign b_s[1075916:1074408] = s_w_712;
assign b_c[1077425:1075917] = c_w_713;assign b_s[1077425:1075917] = s_w_713;
assign b_c[1078934:1077426] = c_w_714;assign b_s[1078934:1077426] = s_w_714;
assign b_c[1080443:1078935] = c_w_715;assign b_s[1080443:1078935] = s_w_715;
assign b_c[1081952:1080444] = c_w_716;assign b_s[1081952:1080444] = s_w_716;
assign b_c[1083461:1081953] = c_w_717;assign b_s[1083461:1081953] = s_w_717;
assign b_c[1084970:1083462] = c_w_718;assign b_s[1084970:1083462] = s_w_718;
assign b_c[1086479:1084971] = c_w_719;assign b_s[1086479:1084971] = s_w_719;
assign b_c[1087988:1086480] = c_w_720;assign b_s[1087988:1086480] = s_w_720;
assign b_c[1089497:1087989] = c_w_721;assign b_s[1089497:1087989] = s_w_721;
assign b_c[1091006:1089498] = c_w_722;assign b_s[1091006:1089498] = s_w_722;
assign b_c[1092515:1091007] = c_w_723;assign b_s[1092515:1091007] = s_w_723;
assign b_c[1094024:1092516] = c_w_724;assign b_s[1094024:1092516] = s_w_724;
assign b_c[1095533:1094025] = c_w_725;assign b_s[1095533:1094025] = s_w_725;
assign b_c[1097042:1095534] = c_w_726;assign b_s[1097042:1095534] = s_w_726;
assign b_c[1098551:1097043] = c_w_727;assign b_s[1098551:1097043] = s_w_727;
assign b_c[1100060:1098552] = c_w_728;assign b_s[1100060:1098552] = s_w_728;
assign b_c[1101569:1100061] = c_w_729;assign b_s[1101569:1100061] = s_w_729;
assign b_c[1103078:1101570] = c_w_730;assign b_s[1103078:1101570] = s_w_730;
assign b_c[1104587:1103079] = c_w_731;assign b_s[1104587:1103079] = s_w_731;
assign b_c[1106096:1104588] = c_w_732;assign b_s[1106096:1104588] = s_w_732;
assign b_c[1107605:1106097] = c_w_733;assign b_s[1107605:1106097] = s_w_733;
assign b_c[1109114:1107606] = c_w_734;assign b_s[1109114:1107606] = s_w_734;
assign b_c[1110623:1109115] = c_w_735;assign b_s[1110623:1109115] = s_w_735;
assign b_c[1112132:1110624] = c_w_736;assign b_s[1112132:1110624] = s_w_736;
assign b_c[1113641:1112133] = c_w_737;assign b_s[1113641:1112133] = s_w_737;
assign b_c[1115150:1113642] = c_w_738;assign b_s[1115150:1113642] = s_w_738;
assign b_c[1116659:1115151] = c_w_739;assign b_s[1116659:1115151] = s_w_739;
assign b_c[1118168:1116660] = c_w_740;assign b_s[1118168:1116660] = s_w_740;
assign b_c[1119677:1118169] = c_w_741;assign b_s[1119677:1118169] = s_w_741;
assign b_c[1121186:1119678] = c_w_742;assign b_s[1121186:1119678] = s_w_742;
assign b_c[1122695:1121187] = c_w_743;assign b_s[1122695:1121187] = s_w_743;
assign b_c[1124204:1122696] = c_w_744;assign b_s[1124204:1122696] = s_w_744;
assign b_c[1125713:1124205] = c_w_745;assign b_s[1125713:1124205] = s_w_745;
assign b_c[1127222:1125714] = c_w_746;assign b_s[1127222:1125714] = s_w_746;
assign b_c[1128731:1127223] = c_w_747;assign b_s[1128731:1127223] = s_w_747;
assign b_c[1130240:1128732] = c_w_748;assign b_s[1130240:1128732] = s_w_748;
assign b_c[1131749:1130241] = c_w_749;assign b_s[1131749:1130241] = s_w_749;
assign b_c[1133258:1131750] = c_w_750;assign b_s[1133258:1131750] = s_w_750;
assign b_c[1134767:1133259] = c_w_751;assign b_s[1134767:1133259] = s_w_751;
assign b_c[1136276:1134768] = c_w_752;assign b_s[1136276:1134768] = s_w_752;
assign b_c[1137785:1136277] = c_w_753;assign b_s[1137785:1136277] = s_w_753;
assign b_c[1139294:1137786] = c_w_754;assign b_s[1139294:1137786] = s_w_754;
assign b_c[1140803:1139295] = c_w_755;assign b_s[1140803:1139295] = s_w_755;
assign b_c[1142312:1140804] = c_w_756;assign b_s[1142312:1140804] = s_w_756;
assign b_c[1143821:1142313] = c_w_757;assign b_s[1143821:1142313] = s_w_757;
assign b_c[1145330:1143822] = c_w_758;assign b_s[1145330:1143822] = s_w_758;
assign b_c[1146839:1145331] = c_w_759;assign b_s[1146839:1145331] = s_w_759;
assign b_c[1148348:1146840] = c_w_760;assign b_s[1148348:1146840] = s_w_760;
assign b_c[1149857:1148349] = c_w_761;assign b_s[1149857:1148349] = s_w_761;
assign b_c[1151366:1149858] = c_w_762;assign b_s[1151366:1149858] = s_w_762;
assign b_c[1152875:1151367] = c_w_763;assign b_s[1152875:1151367] = s_w_763;
assign b_c[1154384:1152876] = c_w_764;assign b_s[1154384:1152876] = s_w_764;
assign b_c[1155893:1154385] = c_w_765;assign b_s[1155893:1154385] = s_w_765;
assign b_c[1157402:1155894] = c_w_766;assign b_s[1157402:1155894] = s_w_766;
assign b_c[1158911:1157403] = c_w_767;assign b_s[1158911:1157403] = s_w_767;
assign b_c[1160420:1158912] = c_w_768;assign b_s[1160420:1158912] = s_w_768;
assign b_c[1161929:1160421] = c_w_769;assign b_s[1161929:1160421] = s_w_769;
assign b_c[1163438:1161930] = c_w_770;assign b_s[1163438:1161930] = s_w_770;
assign b_c[1164947:1163439] = c_w_771;assign b_s[1164947:1163439] = s_w_771;
assign b_c[1166456:1164948] = c_w_772;assign b_s[1166456:1164948] = s_w_772;
assign b_c[1167965:1166457] = c_w_773;assign b_s[1167965:1166457] = s_w_773;
assign b_c[1169474:1167966] = c_w_774;assign b_s[1169474:1167966] = s_w_774;
assign b_c[1170983:1169475] = c_w_775;assign b_s[1170983:1169475] = s_w_775;
assign b_c[1172492:1170984] = c_w_776;assign b_s[1172492:1170984] = s_w_776;
assign b_c[1174001:1172493] = c_w_777;assign b_s[1174001:1172493] = s_w_777;
assign b_c[1175510:1174002] = c_w_778;assign b_s[1175510:1174002] = s_w_778;
assign b_c[1177019:1175511] = c_w_779;assign b_s[1177019:1175511] = s_w_779;
assign b_c[1178528:1177020] = c_w_780;assign b_s[1178528:1177020] = s_w_780;
assign b_c[1180037:1178529] = c_w_781;assign b_s[1180037:1178529] = s_w_781;
assign b_c[1181546:1180038] = c_w_782;assign b_s[1181546:1180038] = s_w_782;
assign b_c[1183055:1181547] = c_w_783;assign b_s[1183055:1181547] = s_w_783;
assign b_c[1184564:1183056] = c_w_784;assign b_s[1184564:1183056] = s_w_784;
assign b_c[1186073:1184565] = c_w_785;assign b_s[1186073:1184565] = s_w_785;
assign b_c[1187582:1186074] = c_w_786;assign b_s[1187582:1186074] = s_w_786;
assign b_c[1189091:1187583] = c_w_787;assign b_s[1189091:1187583] = s_w_787;
assign b_c[1190600:1189092] = c_w_788;assign b_s[1190600:1189092] = s_w_788;
assign b_c[1192109:1190601] = c_w_789;assign b_s[1192109:1190601] = s_w_789;
assign b_c[1193618:1192110] = c_w_790;assign b_s[1193618:1192110] = s_w_790;
assign b_c[1195127:1193619] = c_w_791;assign b_s[1195127:1193619] = s_w_791;
assign b_c[1196636:1195128] = c_w_792;assign b_s[1196636:1195128] = s_w_792;
assign b_c[1198145:1196637] = c_w_793;assign b_s[1198145:1196637] = s_w_793;
assign b_c[1199654:1198146] = c_w_794;assign b_s[1199654:1198146] = s_w_794;
assign b_c[1201163:1199655] = c_w_795;assign b_s[1201163:1199655] = s_w_795;
assign b_c[1202672:1201164] = c_w_796;assign b_s[1202672:1201164] = s_w_796;
assign b_c[1204181:1202673] = c_w_797;assign b_s[1204181:1202673] = s_w_797;
assign b_c[1205690:1204182] = c_w_798;assign b_s[1205690:1204182] = s_w_798;
assign b_c[1207199:1205691] = c_w_799;assign b_s[1207199:1205691] = s_w_799;
assign b_c[1208708:1207200] = c_w_800;assign b_s[1208708:1207200] = s_w_800;
assign b_c[1210217:1208709] = c_w_801;assign b_s[1210217:1208709] = s_w_801;
assign b_c[1211726:1210218] = c_w_802;assign b_s[1211726:1210218] = s_w_802;
assign b_c[1213235:1211727] = c_w_803;assign b_s[1213235:1211727] = s_w_803;
assign b_c[1214744:1213236] = c_w_804;assign b_s[1214744:1213236] = s_w_804;
assign b_c[1216253:1214745] = c_w_805;assign b_s[1216253:1214745] = s_w_805;
assign b_c[1217762:1216254] = c_w_806;assign b_s[1217762:1216254] = s_w_806;
assign b_c[1219271:1217763] = c_w_807;assign b_s[1219271:1217763] = s_w_807;
assign b_c[1220780:1219272] = c_w_808;assign b_s[1220780:1219272] = s_w_808;
assign b_c[1222289:1220781] = c_w_809;assign b_s[1222289:1220781] = s_w_809;
assign b_c[1223798:1222290] = c_w_810;assign b_s[1223798:1222290] = s_w_810;
assign b_c[1225307:1223799] = c_w_811;assign b_s[1225307:1223799] = s_w_811;
assign b_c[1226816:1225308] = c_w_812;assign b_s[1226816:1225308] = s_w_812;
assign b_c[1228325:1226817] = c_w_813;assign b_s[1228325:1226817] = s_w_813;
assign b_c[1229834:1228326] = c_w_814;assign b_s[1229834:1228326] = s_w_814;
assign b_c[1231343:1229835] = c_w_815;assign b_s[1231343:1229835] = s_w_815;
assign b_c[1232852:1231344] = c_w_816;assign b_s[1232852:1231344] = s_w_816;
assign b_c[1234361:1232853] = c_w_817;assign b_s[1234361:1232853] = s_w_817;
assign b_c[1235870:1234362] = c_w_818;assign b_s[1235870:1234362] = s_w_818;
assign b_c[1237379:1235871] = c_w_819;assign b_s[1237379:1235871] = s_w_819;
assign b_c[1238888:1237380] = c_w_820;assign b_s[1238888:1237380] = s_w_820;
assign b_c[1240397:1238889] = c_w_821;assign b_s[1240397:1238889] = s_w_821;
assign b_c[1241906:1240398] = c_w_822;assign b_s[1241906:1240398] = s_w_822;
assign b_c[1243415:1241907] = c_w_823;assign b_s[1243415:1241907] = s_w_823;
assign b_c[1244924:1243416] = c_w_824;assign b_s[1244924:1243416] = s_w_824;
assign b_c[1246433:1244925] = c_w_825;assign b_s[1246433:1244925] = s_w_825;
assign b_c[1247942:1246434] = c_w_826;assign b_s[1247942:1246434] = s_w_826;
assign b_c[1249451:1247943] = c_w_827;assign b_s[1249451:1247943] = s_w_827;
assign b_c[1250960:1249452] = c_w_828;assign b_s[1250960:1249452] = s_w_828;
assign b_c[1252469:1250961] = c_w_829;assign b_s[1252469:1250961] = s_w_829;
assign b_c[1253978:1252470] = c_w_830;assign b_s[1253978:1252470] = s_w_830;
assign b_c[1255487:1253979] = c_w_831;assign b_s[1255487:1253979] = s_w_831;
assign b_c[1256996:1255488] = c_w_832;assign b_s[1256996:1255488] = s_w_832;
assign b_c[1258505:1256997] = c_w_833;assign b_s[1258505:1256997] = s_w_833;
assign b_c[1260014:1258506] = c_w_834;assign b_s[1260014:1258506] = s_w_834;
assign b_c[1261523:1260015] = c_w_835;assign b_s[1261523:1260015] = s_w_835;
assign b_c[1263032:1261524] = c_w_836;assign b_s[1263032:1261524] = s_w_836;
assign b_c[1264541:1263033] = c_w_837;assign b_s[1264541:1263033] = s_w_837;
assign b_c[1266050:1264542] = c_w_838;assign b_s[1266050:1264542] = s_w_838;
assign b_c[1267559:1266051] = c_w_839;assign b_s[1267559:1266051] = s_w_839;
assign b_c[1269068:1267560] = c_w_840;assign b_s[1269068:1267560] = s_w_840;
assign b_c[1270577:1269069] = c_w_841;assign b_s[1270577:1269069] = s_w_841;
assign b_c[1272086:1270578] = c_w_842;assign b_s[1272086:1270578] = s_w_842;
assign b_c[1273595:1272087] = c_w_843;assign b_s[1273595:1272087] = s_w_843;
assign b_c[1275104:1273596] = c_w_844;assign b_s[1275104:1273596] = s_w_844;
assign b_c[1276613:1275105] = c_w_845;assign b_s[1276613:1275105] = s_w_845;
assign b_c[1278122:1276614] = c_w_846;assign b_s[1278122:1276614] = s_w_846;
assign b_c[1279631:1278123] = c_w_847;assign b_s[1279631:1278123] = s_w_847;
assign b_c[1281140:1279632] = c_w_848;assign b_s[1281140:1279632] = s_w_848;
assign b_c[1282649:1281141] = c_w_849;assign b_s[1282649:1281141] = s_w_849;
assign b_c[1284158:1282650] = c_w_850;assign b_s[1284158:1282650] = s_w_850;
assign b_c[1285667:1284159] = c_w_851;assign b_s[1285667:1284159] = s_w_851;
assign b_c[1287176:1285668] = c_w_852;assign b_s[1287176:1285668] = s_w_852;
assign b_c[1288685:1287177] = c_w_853;assign b_s[1288685:1287177] = s_w_853;
assign b_c[1290194:1288686] = c_w_854;assign b_s[1290194:1288686] = s_w_854;
assign b_c[1291703:1290195] = c_w_855;assign b_s[1291703:1290195] = s_w_855;
assign b_c[1293212:1291704] = c_w_856;assign b_s[1293212:1291704] = s_w_856;
assign b_c[1294721:1293213] = c_w_857;assign b_s[1294721:1293213] = s_w_857;
assign b_c[1296230:1294722] = c_w_858;assign b_s[1296230:1294722] = s_w_858;
assign b_c[1297739:1296231] = c_w_859;assign b_s[1297739:1296231] = s_w_859;
assign b_c[1299248:1297740] = c_w_860;assign b_s[1299248:1297740] = s_w_860;
assign b_c[1300757:1299249] = c_w_861;assign b_s[1300757:1299249] = s_w_861;
assign b_c[1302266:1300758] = c_w_862;assign b_s[1302266:1300758] = s_w_862;
assign b_c[1303775:1302267] = c_w_863;assign b_s[1303775:1302267] = s_w_863;
assign b_c[1305284:1303776] = c_w_864;assign b_s[1305284:1303776] = s_w_864;
assign b_c[1306793:1305285] = c_w_865;assign b_s[1306793:1305285] = s_w_865;
assign b_c[1308302:1306794] = c_w_866;assign b_s[1308302:1306794] = s_w_866;
assign b_c[1309811:1308303] = c_w_867;assign b_s[1309811:1308303] = s_w_867;
assign b_c[1311320:1309812] = c_w_868;assign b_s[1311320:1309812] = s_w_868;
assign b_c[1312829:1311321] = c_w_869;assign b_s[1312829:1311321] = s_w_869;
assign b_c[1314338:1312830] = c_w_870;assign b_s[1314338:1312830] = s_w_870;
assign b_c[1315847:1314339] = c_w_871;assign b_s[1315847:1314339] = s_w_871;
assign b_c[1317356:1315848] = c_w_872;assign b_s[1317356:1315848] = s_w_872;
assign b_c[1318865:1317357] = c_w_873;assign b_s[1318865:1317357] = s_w_873;
assign b_c[1320374:1318866] = c_w_874;assign b_s[1320374:1318866] = s_w_874;
assign b_c[1321883:1320375] = c_w_875;assign b_s[1321883:1320375] = s_w_875;
assign b_c[1323392:1321884] = c_w_876;assign b_s[1323392:1321884] = s_w_876;
assign b_c[1324901:1323393] = c_w_877;assign b_s[1324901:1323393] = s_w_877;
assign b_c[1326410:1324902] = c_w_878;assign b_s[1326410:1324902] = s_w_878;
assign b_c[1327919:1326411] = c_w_879;assign b_s[1327919:1326411] = s_w_879;
assign b_c[1329428:1327920] = c_w_880;assign b_s[1329428:1327920] = s_w_880;
assign b_c[1330937:1329429] = c_w_881;assign b_s[1330937:1329429] = s_w_881;
assign b_c[1332446:1330938] = c_w_882;assign b_s[1332446:1330938] = s_w_882;
assign b_c[1333955:1332447] = c_w_883;assign b_s[1333955:1332447] = s_w_883;
assign b_c[1335464:1333956] = c_w_884;assign b_s[1335464:1333956] = s_w_884;
assign b_c[1336973:1335465] = c_w_885;assign b_s[1336973:1335465] = s_w_885;
assign b_c[1338482:1336974] = c_w_886;assign b_s[1338482:1336974] = s_w_886;
assign b_c[1339991:1338483] = c_w_887;assign b_s[1339991:1338483] = s_w_887;
assign b_c[1341500:1339992] = c_w_888;assign b_s[1341500:1339992] = s_w_888;
assign b_c[1343009:1341501] = c_w_889;assign b_s[1343009:1341501] = s_w_889;
assign b_c[1344518:1343010] = c_w_890;assign b_s[1344518:1343010] = s_w_890;
assign b_c[1346027:1344519] = c_w_891;assign b_s[1346027:1344519] = s_w_891;
assign b_c[1347536:1346028] = c_w_892;assign b_s[1347536:1346028] = s_w_892;
assign b_c[1349045:1347537] = c_w_893;assign b_s[1349045:1347537] = s_w_893;
assign b_c[1350554:1349046] = c_w_894;assign b_s[1350554:1349046] = s_w_894;
assign b_c[1352063:1350555] = c_w_895;assign b_s[1352063:1350555] = s_w_895;
assign b_c[1353572:1352064] = c_w_896;assign b_s[1353572:1352064] = s_w_896;
assign b_c[1355081:1353573] = c_w_897;assign b_s[1355081:1353573] = s_w_897;
assign b_c[1356590:1355082] = c_w_898;assign b_s[1356590:1355082] = s_w_898;
assign b_c[1358099:1356591] = c_w_899;assign b_s[1358099:1356591] = s_w_899;
assign b_c[1359608:1358100] = c_w_900;assign b_s[1359608:1358100] = s_w_900;
assign b_c[1361117:1359609] = c_w_901;assign b_s[1361117:1359609] = s_w_901;
assign b_c[1362626:1361118] = c_w_902;assign b_s[1362626:1361118] = s_w_902;
assign b_c[1364135:1362627] = c_w_903;assign b_s[1364135:1362627] = s_w_903;
assign b_c[1365644:1364136] = c_w_904;assign b_s[1365644:1364136] = s_w_904;
assign b_c[1367153:1365645] = c_w_905;assign b_s[1367153:1365645] = s_w_905;
assign b_c[1368662:1367154] = c_w_906;assign b_s[1368662:1367154] = s_w_906;
assign b_c[1370171:1368663] = c_w_907;assign b_s[1370171:1368663] = s_w_907;
assign b_c[1371680:1370172] = c_w_908;assign b_s[1371680:1370172] = s_w_908;
assign b_c[1373189:1371681] = c_w_909;assign b_s[1373189:1371681] = s_w_909;
assign b_c[1374698:1373190] = c_w_910;assign b_s[1374698:1373190] = s_w_910;
assign b_c[1376207:1374699] = c_w_911;assign b_s[1376207:1374699] = s_w_911;
assign b_c[1377716:1376208] = c_w_912;assign b_s[1377716:1376208] = s_w_912;
assign b_c[1379225:1377717] = c_w_913;assign b_s[1379225:1377717] = s_w_913;
assign b_c[1380734:1379226] = c_w_914;assign b_s[1380734:1379226] = s_w_914;
assign b_c[1382243:1380735] = c_w_915;assign b_s[1382243:1380735] = s_w_915;
assign b_c[1383752:1382244] = c_w_916;assign b_s[1383752:1382244] = s_w_916;
assign b_c[1385261:1383753] = c_w_917;assign b_s[1385261:1383753] = s_w_917;
assign b_c[1386770:1385262] = c_w_918;assign b_s[1386770:1385262] = s_w_918;
assign b_c[1388279:1386771] = c_w_919;assign b_s[1388279:1386771] = s_w_919;
assign b_c[1389788:1388280] = c_w_920;assign b_s[1389788:1388280] = s_w_920;
assign b_c[1391297:1389789] = c_w_921;assign b_s[1391297:1389789] = s_w_921;
assign b_c[1392806:1391298] = c_w_922;assign b_s[1392806:1391298] = s_w_922;
assign b_c[1394315:1392807] = c_w_923;assign b_s[1394315:1392807] = s_w_923;
assign b_c[1395824:1394316] = c_w_924;assign b_s[1395824:1394316] = s_w_924;
assign b_c[1397333:1395825] = c_w_925;assign b_s[1397333:1395825] = s_w_925;
assign b_c[1398842:1397334] = c_w_926;assign b_s[1398842:1397334] = s_w_926;
assign b_c[1400351:1398843] = c_w_927;assign b_s[1400351:1398843] = s_w_927;
assign b_c[1401860:1400352] = c_w_928;assign b_s[1401860:1400352] = s_w_928;
assign b_c[1403369:1401861] = c_w_929;assign b_s[1403369:1401861] = s_w_929;
assign b_c[1404878:1403370] = c_w_930;assign b_s[1404878:1403370] = s_w_930;
assign b_c[1406387:1404879] = c_w_931;assign b_s[1406387:1404879] = s_w_931;
assign b_c[1407896:1406388] = c_w_932;assign b_s[1407896:1406388] = s_w_932;
assign b_c[1409405:1407897] = c_w_933;assign b_s[1409405:1407897] = s_w_933;
assign b_c[1410914:1409406] = c_w_934;assign b_s[1410914:1409406] = s_w_934;
assign b_c[1412423:1410915] = c_w_935;assign b_s[1412423:1410915] = s_w_935;
assign b_c[1413932:1412424] = c_w_936;assign b_s[1413932:1412424] = s_w_936;
assign b_c[1415441:1413933] = c_w_937;assign b_s[1415441:1413933] = s_w_937;
assign b_c[1416950:1415442] = c_w_938;assign b_s[1416950:1415442] = s_w_938;
assign b_c[1418459:1416951] = c_w_939;assign b_s[1418459:1416951] = s_w_939;
assign b_c[1419968:1418460] = c_w_940;assign b_s[1419968:1418460] = s_w_940;
assign b_c[1421477:1419969] = c_w_941;assign b_s[1421477:1419969] = s_w_941;
assign b_c[1422986:1421478] = c_w_942;assign b_s[1422986:1421478] = s_w_942;
assign b_c[1424495:1422987] = c_w_943;assign b_s[1424495:1422987] = s_w_943;
assign b_c[1426004:1424496] = c_w_944;assign b_s[1426004:1424496] = s_w_944;
assign b_c[1427513:1426005] = c_w_945;assign b_s[1427513:1426005] = s_w_945;
assign b_c[1429022:1427514] = c_w_946;assign b_s[1429022:1427514] = s_w_946;
assign b_c[1430531:1429023] = c_w_947;assign b_s[1430531:1429023] = s_w_947;
assign b_c[1432040:1430532] = c_w_948;assign b_s[1432040:1430532] = s_w_948;
assign b_c[1433549:1432041] = c_w_949;assign b_s[1433549:1432041] = s_w_949;
assign b_c[1435058:1433550] = c_w_950;assign b_s[1435058:1433550] = s_w_950;
assign b_c[1436567:1435059] = c_w_951;assign b_s[1436567:1435059] = s_w_951;
assign b_c[1438076:1436568] = c_w_952;assign b_s[1438076:1436568] = s_w_952;
assign b_c[1439585:1438077] = c_w_953;assign b_s[1439585:1438077] = s_w_953;
assign b_c[1441094:1439586] = c_w_954;assign b_s[1441094:1439586] = s_w_954;
assign b_c[1442603:1441095] = c_w_955;assign b_s[1442603:1441095] = s_w_955;
assign b_c[1444112:1442604] = c_w_956;assign b_s[1444112:1442604] = s_w_956;
assign b_c[1445621:1444113] = c_w_957;assign b_s[1445621:1444113] = s_w_957;
assign b_c[1447130:1445622] = c_w_958;assign b_s[1447130:1445622] = s_w_958;
assign b_c[1448639:1447131] = c_w_959;assign b_s[1448639:1447131] = s_w_959;
assign b_c[1450148:1448640] = c_w_960;assign b_s[1450148:1448640] = s_w_960;
assign b_c[1451657:1450149] = c_w_961;assign b_s[1451657:1450149] = s_w_961;
assign b_c[1453166:1451658] = c_w_962;assign b_s[1453166:1451658] = s_w_962;
assign b_c[1454675:1453167] = c_w_963;assign b_s[1454675:1453167] = s_w_963;
assign b_c[1456184:1454676] = c_w_964;assign b_s[1456184:1454676] = s_w_964;
assign b_c[1457693:1456185] = c_w_965;assign b_s[1457693:1456185] = s_w_965;
assign b_c[1459202:1457694] = c_w_966;assign b_s[1459202:1457694] = s_w_966;
assign b_c[1460711:1459203] = c_w_967;assign b_s[1460711:1459203] = s_w_967;
assign b_c[1462220:1460712] = c_w_968;assign b_s[1462220:1460712] = s_w_968;
assign b_c[1463729:1462221] = c_w_969;assign b_s[1463729:1462221] = s_w_969;
assign b_c[1465238:1463730] = c_w_970;assign b_s[1465238:1463730] = s_w_970;
assign b_c[1466747:1465239] = c_w_971;assign b_s[1466747:1465239] = s_w_971;
assign b_c[1468256:1466748] = c_w_972;assign b_s[1468256:1466748] = s_w_972;
assign b_c[1469765:1468257] = c_w_973;assign b_s[1469765:1468257] = s_w_973;
assign b_c[1471274:1469766] = c_w_974;assign b_s[1471274:1469766] = s_w_974;
assign b_c[1472783:1471275] = c_w_975;assign b_s[1472783:1471275] = s_w_975;
assign b_c[1474292:1472784] = c_w_976;assign b_s[1474292:1472784] = s_w_976;
assign b_c[1475801:1474293] = c_w_977;assign b_s[1475801:1474293] = s_w_977;
assign b_c[1477310:1475802] = c_w_978;assign b_s[1477310:1475802] = s_w_978;
assign b_c[1478819:1477311] = c_w_979;assign b_s[1478819:1477311] = s_w_979;
assign b_c[1480328:1478820] = c_w_980;assign b_s[1480328:1478820] = s_w_980;
assign b_c[1481837:1480329] = c_w_981;assign b_s[1481837:1480329] = s_w_981;
assign b_c[1483346:1481838] = c_w_982;assign b_s[1483346:1481838] = s_w_982;
assign b_c[1484855:1483347] = c_w_983;assign b_s[1484855:1483347] = s_w_983;
assign b_c[1486364:1484856] = c_w_984;assign b_s[1486364:1484856] = s_w_984;
assign b_c[1487873:1486365] = c_w_985;assign b_s[1487873:1486365] = s_w_985;
assign b_c[1489382:1487874] = c_w_986;assign b_s[1489382:1487874] = s_w_986;
assign b_c[1490891:1489383] = c_w_987;assign b_s[1490891:1489383] = s_w_987;
assign b_c[1492400:1490892] = c_w_988;assign b_s[1492400:1490892] = s_w_988;
assign b_c[1493909:1492401] = c_w_989;assign b_s[1493909:1492401] = s_w_989;
assign b_c[1495418:1493910] = c_w_990;assign b_s[1495418:1493910] = s_w_990;
assign b_c[1496927:1495419] = c_w_991;assign b_s[1496927:1495419] = s_w_991;
assign b_c[1498436:1496928] = c_w_992;assign b_s[1498436:1496928] = s_w_992;
assign b_c[1499945:1498437] = c_w_993;assign b_s[1499945:1498437] = s_w_993;
assign b_c[1501454:1499946] = c_w_994;assign b_s[1501454:1499946] = s_w_994;
assign b_c[1502963:1501455] = c_w_995;assign b_s[1502963:1501455] = s_w_995;
assign b_c[1504472:1502964] = c_w_996;assign b_s[1504472:1502964] = s_w_996;
assign b_c[1505981:1504473] = c_w_997;assign b_s[1505981:1504473] = s_w_997;
assign b_c[1507490:1505982] = c_w_998;assign b_s[1507490:1505982] = s_w_998;
assign b_c[1508999:1507491] = c_w_999;assign b_s[1508999:1507491] = s_w_999;
assign b_c[1510508:1509000] = c_w_1000;assign b_s[1510508:1509000] = s_w_1000;
assign b_c[1512017:1510509] = c_w_1001;assign b_s[1512017:1510509] = s_w_1001;
assign b_c[1513526:1512018] = c_w_1002;assign b_s[1513526:1512018] = s_w_1002;
assign b_c[1515035:1513527] = c_w_1003;assign b_s[1515035:1513527] = s_w_1003;
assign b_c[1516544:1515036] = c_w_1004;assign b_s[1516544:1515036] = s_w_1004;
assign b_c[1518053:1516545] = c_w_1005;assign b_s[1518053:1516545] = s_w_1005;
assign b_c[1519562:1518054] = c_w_1006;assign b_s[1519562:1518054] = s_w_1006;
assign b_c[1521071:1519563] = c_w_1007;assign b_s[1521071:1519563] = s_w_1007;
assign b_c[1522580:1521072] = c_w_1008;assign b_s[1522580:1521072] = s_w_1008;
assign b_c[1524089:1522581] = c_w_1009;assign b_s[1524089:1522581] = s_w_1009;
assign b_c[1525598:1524090] = c_w_1010;assign b_s[1525598:1524090] = s_w_1010;
assign b_c[1527107:1525599] = c_w_1011;assign b_s[1527107:1525599] = s_w_1011;
assign b_c[1528616:1527108] = c_w_1012;assign b_s[1528616:1527108] = s_w_1012;
assign b_c[1530125:1528617] = c_w_1013;assign b_s[1530125:1528617] = s_w_1013;
assign b_c[1531634:1530126] = c_w_1014;assign b_s[1531634:1530126] = s_w_1014;
assign b_c[1533143:1531635] = c_w_1015;assign b_s[1533143:1531635] = s_w_1015;
assign b_c[1534652:1533144] = c_w_1016;assign b_s[1534652:1533144] = s_w_1016;
assign b_c[1536161:1534653] = c_w_1017;assign b_s[1536161:1534653] = s_w_1017;
assign b_c[1537670:1536162] = c_w_1018;assign b_s[1537670:1536162] = s_w_1018;
assign b_c[1539179:1537671] = c_w_1019;assign b_s[1539179:1537671] = s_w_1019;
assign b_c[1540688:1539180] = c_w_1020;assign b_s[1540688:1539180] = s_w_1020;
assign b_c[1542197:1540689] = c_w_1021;assign b_s[1542197:1540689] = s_w_1021;
assign b_c[1543706:1542198] = c_w_1022;assign b_s[1543706:1542198] = s_w_1022;
assign b_c[1545215:1543707] = c_w_1023;assign b_s[1545215:1543707] = s_w_1023;
assign b_c[1546724:1545216] = c_w_1024;assign b_s[1546724:1545216] = s_w_1024;
assign b_c[1548233:1546725] = c_w_1025;assign b_s[1548233:1546725] = s_w_1025;
assign b_c[1549742:1548234] = c_w_1026;assign b_s[1549742:1548234] = s_w_1026;
assign b_c[1551251:1549743] = c_w_1027;assign b_s[1551251:1549743] = s_w_1027;
assign b_c[1552760:1551252] = c_w_1028;assign b_s[1552760:1551252] = s_w_1028;
assign b_c[1554269:1552761] = c_w_1029;assign b_s[1554269:1552761] = s_w_1029;
assign b_c[1555778:1554270] = c_w_1030;assign b_s[1555778:1554270] = s_w_1030;
assign b_c[1557287:1555779] = c_w_1031;assign b_s[1557287:1555779] = s_w_1031;
assign b_c[1558796:1557288] = c_w_1032;assign b_s[1558796:1557288] = s_w_1032;
assign b_c[1560305:1558797] = c_w_1033;assign b_s[1560305:1558797] = s_w_1033;
assign b_c[1561814:1560306] = c_w_1034;assign b_s[1561814:1560306] = s_w_1034;
assign b_c[1563323:1561815] = c_w_1035;assign b_s[1563323:1561815] = s_w_1035;
assign b_c[1564832:1563324] = c_w_1036;assign b_s[1564832:1563324] = s_w_1036;
assign b_c[1566341:1564833] = c_w_1037;assign b_s[1566341:1564833] = s_w_1037;
assign b_c[1567850:1566342] = c_w_1038;assign b_s[1567850:1566342] = s_w_1038;
assign b_c[1569359:1567851] = c_w_1039;assign b_s[1569359:1567851] = s_w_1039;
assign b_c[1570868:1569360] = c_w_1040;assign b_s[1570868:1569360] = s_w_1040;
assign b_c[1572377:1570869] = c_w_1041;assign b_s[1572377:1570869] = s_w_1041;
assign b_c[1573886:1572378] = c_w_1042;assign b_s[1573886:1572378] = s_w_1042;
assign b_c[1575395:1573887] = c_w_1043;assign b_s[1575395:1573887] = s_w_1043;
assign b_c[1576904:1575396] = c_w_1044;assign b_s[1576904:1575396] = s_w_1044;
assign b_c[1578413:1576905] = c_w_1045;assign b_s[1578413:1576905] = s_w_1045;
assign b_c[1579922:1578414] = c_w_1046;assign b_s[1579922:1578414] = s_w_1046;
assign b_c[1581431:1579923] = c_w_1047;assign b_s[1581431:1579923] = s_w_1047;
assign b_c[1582940:1581432] = c_w_1048;assign b_s[1582940:1581432] = s_w_1048;
assign b_c[1584449:1582941] = c_w_1049;assign b_s[1584449:1582941] = s_w_1049;
assign b_c[1585958:1584450] = c_w_1050;assign b_s[1585958:1584450] = s_w_1050;
assign b_c[1587467:1585959] = c_w_1051;assign b_s[1587467:1585959] = s_w_1051;
assign b_c[1588976:1587468] = c_w_1052;assign b_s[1588976:1587468] = s_w_1052;
assign b_c[1590485:1588977] = c_w_1053;assign b_s[1590485:1588977] = s_w_1053;
assign b_c[1591994:1590486] = c_w_1054;assign b_s[1591994:1590486] = s_w_1054;
assign b_c[1593503:1591995] = c_w_1055;assign b_s[1593503:1591995] = s_w_1055;
assign b_c[1595012:1593504] = c_w_1056;assign b_s[1595012:1593504] = s_w_1056;
assign b_c[1596521:1595013] = c_w_1057;assign b_s[1596521:1595013] = s_w_1057;
assign b_c[1598030:1596522] = c_w_1058;assign b_s[1598030:1596522] = s_w_1058;
assign b_c[1599539:1598031] = c_w_1059;assign b_s[1599539:1598031] = s_w_1059;
assign b_c[1601048:1599540] = c_w_1060;assign b_s[1601048:1599540] = s_w_1060;
assign b_c[1602557:1601049] = c_w_1061;assign b_s[1602557:1601049] = s_w_1061;
assign b_c[1604066:1602558] = c_w_1062;assign b_s[1604066:1602558] = s_w_1062;
assign b_c[1605575:1604067] = c_w_1063;assign b_s[1605575:1604067] = s_w_1063;
assign b_c[1607084:1605576] = c_w_1064;assign b_s[1607084:1605576] = s_w_1064;
assign b_c[1608593:1607085] = c_w_1065;assign b_s[1608593:1607085] = s_w_1065;
assign b_c[1610102:1608594] = c_w_1066;assign b_s[1610102:1608594] = s_w_1066;
assign b_c[1611611:1610103] = c_w_1067;assign b_s[1611611:1610103] = s_w_1067;
assign b_c[1613120:1611612] = c_w_1068;assign b_s[1613120:1611612] = s_w_1068;
assign b_c[1614629:1613121] = c_w_1069;assign b_s[1614629:1613121] = s_w_1069;
assign b_c[1616138:1614630] = c_w_1070;assign b_s[1616138:1614630] = s_w_1070;
assign b_c[1617647:1616139] = c_w_1071;assign b_s[1617647:1616139] = s_w_1071;
assign b_c[1619156:1617648] = c_w_1072;assign b_s[1619156:1617648] = s_w_1072;
assign b_c[1620665:1619157] = c_w_1073;assign b_s[1620665:1619157] = s_w_1073;
assign b_c[1622174:1620666] = c_w_1074;assign b_s[1622174:1620666] = s_w_1074;
assign b_c[1623683:1622175] = c_w_1075;assign b_s[1623683:1622175] = s_w_1075;
assign b_c[1625192:1623684] = c_w_1076;assign b_s[1625192:1623684] = s_w_1076;
assign b_c[1626701:1625193] = c_w_1077;assign b_s[1626701:1625193] = s_w_1077;
assign b_c[1628210:1626702] = c_w_1078;assign b_s[1628210:1626702] = s_w_1078;
assign b_c[1629719:1628211] = c_w_1079;assign b_s[1629719:1628211] = s_w_1079;
assign b_c[1631228:1629720] = c_w_1080;assign b_s[1631228:1629720] = s_w_1080;
assign b_c[1632737:1631229] = c_w_1081;assign b_s[1632737:1631229] = s_w_1081;
assign b_c[1634246:1632738] = c_w_1082;assign b_s[1634246:1632738] = s_w_1082;
assign b_c[1635755:1634247] = c_w_1083;assign b_s[1635755:1634247] = s_w_1083;
assign b_c[1637264:1635756] = c_w_1084;assign b_s[1637264:1635756] = s_w_1084;
assign b_c[1638773:1637265] = c_w_1085;assign b_s[1638773:1637265] = s_w_1085;
assign b_c[1640282:1638774] = c_w_1086;assign b_s[1640282:1638774] = s_w_1086;
assign b_c[1641791:1640283] = c_w_1087;assign b_s[1641791:1640283] = s_w_1087;
assign b_c[1643300:1641792] = c_w_1088;assign b_s[1643300:1641792] = s_w_1088;
assign b_c[1644809:1643301] = c_w_1089;assign b_s[1644809:1643301] = s_w_1089;
assign b_c[1646318:1644810] = c_w_1090;assign b_s[1646318:1644810] = s_w_1090;
assign b_c[1647827:1646319] = c_w_1091;assign b_s[1647827:1646319] = s_w_1091;
assign b_c[1649336:1647828] = c_w_1092;assign b_s[1649336:1647828] = s_w_1092;
assign b_c[1650845:1649337] = c_w_1093;assign b_s[1650845:1649337] = s_w_1093;
assign b_c[1652354:1650846] = c_w_1094;assign b_s[1652354:1650846] = s_w_1094;
assign b_c[1653863:1652355] = c_w_1095;assign b_s[1653863:1652355] = s_w_1095;
assign b_c[1655372:1653864] = c_w_1096;assign b_s[1655372:1653864] = s_w_1096;
assign b_c[1656881:1655373] = c_w_1097;assign b_s[1656881:1655373] = s_w_1097;
assign b_c[1658390:1656882] = c_w_1098;assign b_s[1658390:1656882] = s_w_1098;
assign b_c[1659899:1658391] = c_w_1099;assign b_s[1659899:1658391] = s_w_1099;
assign b_c[1661408:1659900] = c_w_1100;assign b_s[1661408:1659900] = s_w_1100;
assign b_c[1662917:1661409] = c_w_1101;assign b_s[1662917:1661409] = s_w_1101;
assign b_c[1664426:1662918] = c_w_1102;assign b_s[1664426:1662918] = s_w_1102;
assign b_c[1665935:1664427] = c_w_1103;assign b_s[1665935:1664427] = s_w_1103;
assign b_c[1667444:1665936] = c_w_1104;assign b_s[1667444:1665936] = s_w_1104;
assign b_c[1668953:1667445] = c_w_1105;assign b_s[1668953:1667445] = s_w_1105;
assign b_c[1670462:1668954] = c_w_1106;assign b_s[1670462:1668954] = s_w_1106;
assign b_c[1671971:1670463] = c_w_1107;assign b_s[1671971:1670463] = s_w_1107;
assign b_c[1673480:1671972] = c_w_1108;assign b_s[1673480:1671972] = s_w_1108;
assign b_c[1674989:1673481] = c_w_1109;assign b_s[1674989:1673481] = s_w_1109;
assign b_c[1676498:1674990] = c_w_1110;assign b_s[1676498:1674990] = s_w_1110;
assign b_c[1678007:1676499] = c_w_1111;assign b_s[1678007:1676499] = s_w_1111;
assign b_c[1679516:1678008] = c_w_1112;assign b_s[1679516:1678008] = s_w_1112;
assign b_c[1681025:1679517] = c_w_1113;assign b_s[1681025:1679517] = s_w_1113;
assign b_c[1682534:1681026] = c_w_1114;assign b_s[1682534:1681026] = s_w_1114;
assign b_c[1684043:1682535] = c_w_1115;assign b_s[1684043:1682535] = s_w_1115;
assign b_c[1685552:1684044] = c_w_1116;assign b_s[1685552:1684044] = s_w_1116;
assign b_c[1687061:1685553] = c_w_1117;assign b_s[1687061:1685553] = s_w_1117;
assign b_c[1688570:1687062] = c_w_1118;assign b_s[1688570:1687062] = s_w_1118;
assign b_c[1690079:1688571] = c_w_1119;assign b_s[1690079:1688571] = s_w_1119;
assign b_c[1691588:1690080] = c_w_1120;assign b_s[1691588:1690080] = s_w_1120;
assign b_c[1693097:1691589] = c_w_1121;assign b_s[1693097:1691589] = s_w_1121;
assign b_c[1694606:1693098] = c_w_1122;assign b_s[1694606:1693098] = s_w_1122;
assign b_c[1696115:1694607] = c_w_1123;assign b_s[1696115:1694607] = s_w_1123;
assign b_c[1697624:1696116] = c_w_1124;assign b_s[1697624:1696116] = s_w_1124;
assign b_c[1699133:1697625] = c_w_1125;assign b_s[1699133:1697625] = s_w_1125;
assign b_c[1700642:1699134] = c_w_1126;assign b_s[1700642:1699134] = s_w_1126;
assign b_c[1702151:1700643] = c_w_1127;assign b_s[1702151:1700643] = s_w_1127;
assign b_c[1703660:1702152] = c_w_1128;assign b_s[1703660:1702152] = s_w_1128;
assign b_c[1705169:1703661] = c_w_1129;assign b_s[1705169:1703661] = s_w_1129;
assign b_c[1706678:1705170] = c_w_1130;assign b_s[1706678:1705170] = s_w_1130;
assign b_c[1708187:1706679] = c_w_1131;assign b_s[1708187:1706679] = s_w_1131;
assign b_c[1709696:1708188] = c_w_1132;assign b_s[1709696:1708188] = s_w_1132;
assign b_c[1711205:1709697] = c_w_1133;assign b_s[1711205:1709697] = s_w_1133;
assign b_c[1712714:1711206] = c_w_1134;assign b_s[1712714:1711206] = s_w_1134;
assign b_c[1714223:1712715] = c_w_1135;assign b_s[1714223:1712715] = s_w_1135;
assign b_c[1715732:1714224] = c_w_1136;assign b_s[1715732:1714224] = s_w_1136;
assign b_c[1717241:1715733] = c_w_1137;assign b_s[1717241:1715733] = s_w_1137;
assign b_c[1718750:1717242] = c_w_1138;assign b_s[1718750:1717242] = s_w_1138;
assign b_c[1720259:1718751] = c_w_1139;assign b_s[1720259:1718751] = s_w_1139;
assign b_c[1721768:1720260] = c_w_1140;assign b_s[1721768:1720260] = s_w_1140;
assign b_c[1723277:1721769] = c_w_1141;assign b_s[1723277:1721769] = s_w_1141;
assign b_c[1724786:1723278] = c_w_1142;assign b_s[1724786:1723278] = s_w_1142;
assign b_c[1726295:1724787] = c_w_1143;assign b_s[1726295:1724787] = s_w_1143;
assign b_c[1727804:1726296] = c_w_1144;assign b_s[1727804:1726296] = s_w_1144;
assign b_c[1729313:1727805] = c_w_1145;assign b_s[1729313:1727805] = s_w_1145;
assign b_c[1730822:1729314] = c_w_1146;assign b_s[1730822:1729314] = s_w_1146;
assign b_c[1732331:1730823] = c_w_1147;assign b_s[1732331:1730823] = s_w_1147;
assign b_c[1733840:1732332] = c_w_1148;assign b_s[1733840:1732332] = s_w_1148;
assign b_c[1735349:1733841] = c_w_1149;assign b_s[1735349:1733841] = s_w_1149;
assign b_c[1736858:1735350] = c_w_1150;assign b_s[1736858:1735350] = s_w_1150;
assign b_c[1738367:1736859] = c_w_1151;assign b_s[1738367:1736859] = s_w_1151;
assign b_c[1739876:1738368] = c_w_1152;assign b_s[1739876:1738368] = s_w_1152;
assign b_c[1741385:1739877] = c_w_1153;assign b_s[1741385:1739877] = s_w_1153;
assign b_c[1742894:1741386] = c_w_1154;assign b_s[1742894:1741386] = s_w_1154;
assign b_c[1744403:1742895] = c_w_1155;assign b_s[1744403:1742895] = s_w_1155;
assign b_c[1745912:1744404] = c_w_1156;assign b_s[1745912:1744404] = s_w_1156;
assign b_c[1747421:1745913] = c_w_1157;assign b_s[1747421:1745913] = s_w_1157;
assign b_c[1748930:1747422] = c_w_1158;assign b_s[1748930:1747422] = s_w_1158;
assign b_c[1750439:1748931] = c_w_1159;assign b_s[1750439:1748931] = s_w_1159;
assign b_c[1751948:1750440] = c_w_1160;assign b_s[1751948:1750440] = s_w_1160;
assign b_c[1753457:1751949] = c_w_1161;assign b_s[1753457:1751949] = s_w_1161;
assign b_c[1754966:1753458] = c_w_1162;assign b_s[1754966:1753458] = s_w_1162;
assign b_c[1756475:1754967] = c_w_1163;assign b_s[1756475:1754967] = s_w_1163;
assign b_c[1757984:1756476] = c_w_1164;assign b_s[1757984:1756476] = s_w_1164;
assign b_c[1759493:1757985] = c_w_1165;assign b_s[1759493:1757985] = s_w_1165;
assign b_c[1761002:1759494] = c_w_1166;assign b_s[1761002:1759494] = s_w_1166;
assign b_c[1762511:1761003] = c_w_1167;assign b_s[1762511:1761003] = s_w_1167;
assign b_c[1764020:1762512] = c_w_1168;assign b_s[1764020:1762512] = s_w_1168;
assign b_c[1765529:1764021] = c_w_1169;assign b_s[1765529:1764021] = s_w_1169;
assign b_c[1767038:1765530] = c_w_1170;assign b_s[1767038:1765530] = s_w_1170;
assign b_c[1768547:1767039] = c_w_1171;assign b_s[1768547:1767039] = s_w_1171;
assign b_c[1770056:1768548] = c_w_1172;assign b_s[1770056:1768548] = s_w_1172;
assign b_c[1771565:1770057] = c_w_1173;assign b_s[1771565:1770057] = s_w_1173;
assign b_c[1773074:1771566] = c_w_1174;assign b_s[1773074:1771566] = s_w_1174;
assign b_c[1774583:1773075] = c_w_1175;assign b_s[1774583:1773075] = s_w_1175;
assign b_c[1776092:1774584] = c_w_1176;assign b_s[1776092:1774584] = s_w_1176;
assign b_c[1777601:1776093] = c_w_1177;assign b_s[1777601:1776093] = s_w_1177;
assign b_c[1779110:1777602] = c_w_1178;assign b_s[1779110:1777602] = s_w_1178;
assign b_c[1780619:1779111] = c_w_1179;assign b_s[1780619:1779111] = s_w_1179;
assign b_c[1782128:1780620] = c_w_1180;assign b_s[1782128:1780620] = s_w_1180;
assign b_c[1783637:1782129] = c_w_1181;assign b_s[1783637:1782129] = s_w_1181;
assign b_c[1785146:1783638] = c_w_1182;assign b_s[1785146:1783638] = s_w_1182;
assign b_c[1786655:1785147] = c_w_1183;assign b_s[1786655:1785147] = s_w_1183;
assign b_c[1788164:1786656] = c_w_1184;assign b_s[1788164:1786656] = s_w_1184;
assign b_c[1789673:1788165] = c_w_1185;assign b_s[1789673:1788165] = s_w_1185;
assign b_c[1791182:1789674] = c_w_1186;assign b_s[1791182:1789674] = s_w_1186;
assign b_c[1792691:1791183] = c_w_1187;assign b_s[1792691:1791183] = s_w_1187;
assign b_c[1794200:1792692] = c_w_1188;assign b_s[1794200:1792692] = s_w_1188;
assign b_c[1795709:1794201] = c_w_1189;assign b_s[1795709:1794201] = s_w_1189;
assign b_c[1797218:1795710] = c_w_1190;assign b_s[1797218:1795710] = s_w_1190;
assign b_c[1798727:1797219] = c_w_1191;assign b_s[1798727:1797219] = s_w_1191;
assign b_c[1800236:1798728] = c_w_1192;assign b_s[1800236:1798728] = s_w_1192;
assign b_c[1801745:1800237] = c_w_1193;assign b_s[1801745:1800237] = s_w_1193;
assign b_c[1803254:1801746] = c_w_1194;assign b_s[1803254:1801746] = s_w_1194;
assign b_c[1804763:1803255] = c_w_1195;assign b_s[1804763:1803255] = s_w_1195;
assign b_c[1806272:1804764] = c_w_1196;assign b_s[1806272:1804764] = s_w_1196;
assign b_c[1807781:1806273] = c_w_1197;assign b_s[1807781:1806273] = s_w_1197;
assign b_c[1809290:1807782] = c_w_1198;assign b_s[1809290:1807782] = s_w_1198;
assign b_c[1810799:1809291] = c_w_1199;assign b_s[1810799:1809291] = s_w_1199;
assign b_c[1812308:1810800] = c_w_1200;assign b_s[1812308:1810800] = s_w_1200;
assign b_c[1813817:1812309] = c_w_1201;assign b_s[1813817:1812309] = s_w_1201;
assign b_c[1815326:1813818] = c_w_1202;assign b_s[1815326:1813818] = s_w_1202;
assign b_c[1816835:1815327] = c_w_1203;assign b_s[1816835:1815327] = s_w_1203;
assign b_c[1818344:1816836] = c_w_1204;assign b_s[1818344:1816836] = s_w_1204;
assign b_c[1819853:1818345] = c_w_1205;assign b_s[1819853:1818345] = s_w_1205;
assign b_c[1821362:1819854] = c_w_1206;assign b_s[1821362:1819854] = s_w_1206;
assign b_c[1822871:1821363] = c_w_1207;assign b_s[1822871:1821363] = s_w_1207;
assign b_c[1824380:1822872] = c_w_1208;assign b_s[1824380:1822872] = s_w_1208;
assign b_c[1825889:1824381] = c_w_1209;assign b_s[1825889:1824381] = s_w_1209;
assign b_c[1827398:1825890] = c_w_1210;assign b_s[1827398:1825890] = s_w_1210;
assign b_c[1828907:1827399] = c_w_1211;assign b_s[1828907:1827399] = s_w_1211;
assign b_c[1830416:1828908] = c_w_1212;assign b_s[1830416:1828908] = s_w_1212;
assign b_c[1831925:1830417] = c_w_1213;assign b_s[1831925:1830417] = s_w_1213;
assign b_c[1833434:1831926] = c_w_1214;assign b_s[1833434:1831926] = s_w_1214;
assign b_c[1834943:1833435] = c_w_1215;assign b_s[1834943:1833435] = s_w_1215;
assign b_c[1836452:1834944] = c_w_1216;assign b_s[1836452:1834944] = s_w_1216;
assign b_c[1837961:1836453] = c_w_1217;assign b_s[1837961:1836453] = s_w_1217;
assign b_c[1839470:1837962] = c_w_1218;assign b_s[1839470:1837962] = s_w_1218;
assign b_c[1840979:1839471] = c_w_1219;assign b_s[1840979:1839471] = s_w_1219;
assign b_c[1842488:1840980] = c_w_1220;assign b_s[1842488:1840980] = s_w_1220;
assign b_c[1843997:1842489] = c_w_1221;assign b_s[1843997:1842489] = s_w_1221;
assign b_c[1845506:1843998] = c_w_1222;assign b_s[1845506:1843998] = s_w_1222;
assign b_c[1847015:1845507] = c_w_1223;assign b_s[1847015:1845507] = s_w_1223;
assign b_c[1848524:1847016] = c_w_1224;assign b_s[1848524:1847016] = s_w_1224;
assign b_c[1850033:1848525] = c_w_1225;assign b_s[1850033:1848525] = s_w_1225;
assign b_c[1851542:1850034] = c_w_1226;assign b_s[1851542:1850034] = s_w_1226;
assign b_c[1853051:1851543] = c_w_1227;assign b_s[1853051:1851543] = s_w_1227;
assign b_c[1854560:1853052] = c_w_1228;assign b_s[1854560:1853052] = s_w_1228;
assign b_c[1856069:1854561] = c_w_1229;assign b_s[1856069:1854561] = s_w_1229;
assign b_c[1857578:1856070] = c_w_1230;assign b_s[1857578:1856070] = s_w_1230;
assign b_c[1859087:1857579] = c_w_1231;assign b_s[1859087:1857579] = s_w_1231;
assign b_c[1860596:1859088] = c_w_1232;assign b_s[1860596:1859088] = s_w_1232;
assign b_c[1862105:1860597] = c_w_1233;assign b_s[1862105:1860597] = s_w_1233;
assign b_c[1863614:1862106] = c_w_1234;assign b_s[1863614:1862106] = s_w_1234;
assign b_c[1865123:1863615] = c_w_1235;assign b_s[1865123:1863615] = s_w_1235;
assign b_c[1866632:1865124] = c_w_1236;assign b_s[1866632:1865124] = s_w_1236;
assign b_c[1868141:1866633] = c_w_1237;assign b_s[1868141:1866633] = s_w_1237;
assign b_c[1869650:1868142] = c_w_1238;assign b_s[1869650:1868142] = s_w_1238;
assign b_c[1871159:1869651] = c_w_1239;assign b_s[1871159:1869651] = s_w_1239;
assign b_c[1872668:1871160] = c_w_1240;assign b_s[1872668:1871160] = s_w_1240;
assign b_c[1874177:1872669] = c_w_1241;assign b_s[1874177:1872669] = s_w_1241;
assign b_c[1875686:1874178] = c_w_1242;assign b_s[1875686:1874178] = s_w_1242;
assign b_c[1877195:1875687] = c_w_1243;assign b_s[1877195:1875687] = s_w_1243;
assign b_c[1878704:1877196] = c_w_1244;assign b_s[1878704:1877196] = s_w_1244;
assign b_c[1880213:1878705] = c_w_1245;assign b_s[1880213:1878705] = s_w_1245;
assign b_c[1881722:1880214] = c_w_1246;assign b_s[1881722:1880214] = s_w_1246;
assign b_c[1883231:1881723] = c_w_1247;assign b_s[1883231:1881723] = s_w_1247;
assign b_c[1884740:1883232] = c_w_1248;assign b_s[1884740:1883232] = s_w_1248;
assign b_c[1886249:1884741] = c_w_1249;assign b_s[1886249:1884741] = s_w_1249;
assign b_c[1887758:1886250] = c_w_1250;assign b_s[1887758:1886250] = s_w_1250;
assign b_c[1889267:1887759] = c_w_1251;assign b_s[1889267:1887759] = s_w_1251;
assign b_c[1890776:1889268] = c_w_1252;assign b_s[1890776:1889268] = s_w_1252;
assign b_c[1892285:1890777] = c_w_1253;assign b_s[1892285:1890777] = s_w_1253;
assign b_c[1893794:1892286] = c_w_1254;assign b_s[1893794:1892286] = s_w_1254;
assign b_c[1895303:1893795] = c_w_1255;assign b_s[1895303:1893795] = s_w_1255;
assign b_c[1896812:1895304] = c_w_1256;assign b_s[1896812:1895304] = s_w_1256;
assign b_c[1898321:1896813] = c_w_1257;assign b_s[1898321:1896813] = s_w_1257;
assign b_c[1899830:1898322] = c_w_1258;assign b_s[1899830:1898322] = s_w_1258;
assign b_c[1901339:1899831] = c_w_1259;assign b_s[1901339:1899831] = s_w_1259;
assign b_c[1902848:1901340] = c_w_1260;assign b_s[1902848:1901340] = s_w_1260;
assign b_c[1904357:1902849] = c_w_1261;assign b_s[1904357:1902849] = s_w_1261;
assign b_c[1905866:1904358] = c_w_1262;assign b_s[1905866:1904358] = s_w_1262;
assign b_c[1907375:1905867] = c_w_1263;assign b_s[1907375:1905867] = s_w_1263;
assign b_c[1908884:1907376] = c_w_1264;assign b_s[1908884:1907376] = s_w_1264;
assign b_c[1910393:1908885] = c_w_1265;assign b_s[1910393:1908885] = s_w_1265;
assign b_c[1911902:1910394] = c_w_1266;assign b_s[1911902:1910394] = s_w_1266;
assign b_c[1913411:1911903] = c_w_1267;assign b_s[1913411:1911903] = s_w_1267;
assign b_c[1914920:1913412] = c_w_1268;assign b_s[1914920:1913412] = s_w_1268;
assign b_c[1916429:1914921] = c_w_1269;assign b_s[1916429:1914921] = s_w_1269;
assign b_c[1917938:1916430] = c_w_1270;assign b_s[1917938:1916430] = s_w_1270;
assign b_c[1919447:1917939] = c_w_1271;assign b_s[1919447:1917939] = s_w_1271;
assign b_c[1920956:1919448] = c_w_1272;assign b_s[1920956:1919448] = s_w_1272;
assign b_c[1922465:1920957] = c_w_1273;assign b_s[1922465:1920957] = s_w_1273;
assign b_c[1923974:1922466] = c_w_1274;assign b_s[1923974:1922466] = s_w_1274;
assign b_c[1925483:1923975] = c_w_1275;assign b_s[1925483:1923975] = s_w_1275;
assign b_c[1926992:1925484] = c_w_1276;assign b_s[1926992:1925484] = s_w_1276;
assign b_c[1928501:1926993] = c_w_1277;assign b_s[1928501:1926993] = s_w_1277;
assign b_c[1930010:1928502] = c_w_1278;assign b_s[1930010:1928502] = s_w_1278;
assign b_c[1931519:1930011] = c_w_1279;assign b_s[1931519:1930011] = s_w_1279;
assign b_c[1933028:1931520] = c_w_1280;assign b_s[1933028:1931520] = s_w_1280;
assign b_c[1934537:1933029] = c_w_1281;assign b_s[1934537:1933029] = s_w_1281;
assign b_c[1936046:1934538] = c_w_1282;assign b_s[1936046:1934538] = s_w_1282;
assign b_c[1937555:1936047] = c_w_1283;assign b_s[1937555:1936047] = s_w_1283;
assign b_c[1939064:1937556] = c_w_1284;assign b_s[1939064:1937556] = s_w_1284;
assign b_c[1940573:1939065] = c_w_1285;assign b_s[1940573:1939065] = s_w_1285;
assign b_c[1942082:1940574] = c_w_1286;assign b_s[1942082:1940574] = s_w_1286;
assign b_c[1943591:1942083] = c_w_1287;assign b_s[1943591:1942083] = s_w_1287;
assign b_c[1945100:1943592] = c_w_1288;assign b_s[1945100:1943592] = s_w_1288;
assign b_c[1946609:1945101] = c_w_1289;assign b_s[1946609:1945101] = s_w_1289;
assign b_c[1948118:1946610] = c_w_1290;assign b_s[1948118:1946610] = s_w_1290;
assign b_c[1949627:1948119] = c_w_1291;assign b_s[1949627:1948119] = s_w_1291;
assign b_c[1951136:1949628] = c_w_1292;assign b_s[1951136:1949628] = s_w_1292;
assign b_c[1952645:1951137] = c_w_1293;assign b_s[1952645:1951137] = s_w_1293;
assign b_c[1954154:1952646] = c_w_1294;assign b_s[1954154:1952646] = s_w_1294;
assign b_c[1955663:1954155] = c_w_1295;assign b_s[1955663:1954155] = s_w_1295;
assign b_c[1957172:1955664] = c_w_1296;assign b_s[1957172:1955664] = s_w_1296;
assign b_c[1958681:1957173] = c_w_1297;assign b_s[1958681:1957173] = s_w_1297;
assign b_c[1960190:1958682] = c_w_1298;assign b_s[1960190:1958682] = s_w_1298;
assign b_c[1961699:1960191] = c_w_1299;assign b_s[1961699:1960191] = s_w_1299;
assign b_c[1963208:1961700] = c_w_1300;assign b_s[1963208:1961700] = s_w_1300;
assign b_c[1964717:1963209] = c_w_1301;assign b_s[1964717:1963209] = s_w_1301;
assign b_c[1966226:1964718] = c_w_1302;assign b_s[1966226:1964718] = s_w_1302;
assign b_c[1967735:1966227] = c_w_1303;assign b_s[1967735:1966227] = s_w_1303;
assign b_c[1969244:1967736] = c_w_1304;assign b_s[1969244:1967736] = s_w_1304;
assign b_c[1970753:1969245] = c_w_1305;assign b_s[1970753:1969245] = s_w_1305;
assign b_c[1972262:1970754] = c_w_1306;assign b_s[1972262:1970754] = s_w_1306;
assign b_c[1973771:1972263] = c_w_1307;assign b_s[1973771:1972263] = s_w_1307;
assign b_c[1975280:1973772] = c_w_1308;assign b_s[1975280:1973772] = s_w_1308;
assign b_c[1976789:1975281] = c_w_1309;assign b_s[1976789:1975281] = s_w_1309;
assign b_c[1978298:1976790] = c_w_1310;assign b_s[1978298:1976790] = s_w_1310;
assign b_c[1979807:1978299] = c_w_1311;assign b_s[1979807:1978299] = s_w_1311;
assign b_c[1981316:1979808] = c_w_1312;assign b_s[1981316:1979808] = s_w_1312;
assign b_c[1982825:1981317] = c_w_1313;assign b_s[1982825:1981317] = s_w_1313;
assign b_c[1984334:1982826] = c_w_1314;assign b_s[1984334:1982826] = s_w_1314;
assign b_c[1985843:1984335] = c_w_1315;assign b_s[1985843:1984335] = s_w_1315;
assign b_c[1987352:1985844] = c_w_1316;assign b_s[1987352:1985844] = s_w_1316;
assign b_c[1988861:1987353] = c_w_1317;assign b_s[1988861:1987353] = s_w_1317;
assign b_c[1990370:1988862] = c_w_1318;assign b_s[1990370:1988862] = s_w_1318;
assign b_c[1991879:1990371] = c_w_1319;assign b_s[1991879:1990371] = s_w_1319;
assign b_c[1993388:1991880] = c_w_1320;assign b_s[1993388:1991880] = s_w_1320;
assign b_c[1994897:1993389] = c_w_1321;assign b_s[1994897:1993389] = s_w_1321;
assign b_c[1996406:1994898] = c_w_1322;assign b_s[1996406:1994898] = s_w_1322;
assign b_c[1997915:1996407] = c_w_1323;assign b_s[1997915:1996407] = s_w_1323;
assign b_c[1999424:1997916] = c_w_1324;assign b_s[1999424:1997916] = s_w_1324;
assign b_c[2000933:1999425] = c_w_1325;assign b_s[2000933:1999425] = s_w_1325;
assign b_c[2002442:2000934] = c_w_1326;assign b_s[2002442:2000934] = s_w_1326;
assign b_c[2003951:2002443] = c_w_1327;assign b_s[2003951:2002443] = s_w_1327;
assign b_c[2005460:2003952] = c_w_1328;assign b_s[2005460:2003952] = s_w_1328;
assign b_c[2006969:2005461] = c_w_1329;assign b_s[2006969:2005461] = s_w_1329;
assign b_c[2008478:2006970] = c_w_1330;assign b_s[2008478:2006970] = s_w_1330;
assign b_c[2009987:2008479] = c_w_1331;assign b_s[2009987:2008479] = s_w_1331;
assign b_c[2011496:2009988] = c_w_1332;assign b_s[2011496:2009988] = s_w_1332;
assign b_c[2013005:2011497] = c_w_1333;assign b_s[2013005:2011497] = s_w_1333;
assign b_c[2014514:2013006] = c_w_1334;assign b_s[2014514:2013006] = s_w_1334;
assign b_c[2016023:2014515] = c_w_1335;assign b_s[2016023:2014515] = s_w_1335;
assign b_c[2017532:2016024] = c_w_1336;assign b_s[2017532:2016024] = s_w_1336;
assign b_c[2019041:2017533] = c_w_1337;assign b_s[2019041:2017533] = s_w_1337;
assign b_c[2020550:2019042] = c_w_1338;assign b_s[2020550:2019042] = s_w_1338;
assign b_c[2022059:2020551] = c_w_1339;assign b_s[2022059:2020551] = s_w_1339;
assign b_c[2023568:2022060] = c_w_1340;assign b_s[2023568:2022060] = s_w_1340;
assign b_c[2025077:2023569] = c_w_1341;assign b_s[2025077:2023569] = s_w_1341;
assign b_c[2026586:2025078] = c_w_1342;assign b_s[2026586:2025078] = s_w_1342;
assign b_c[2028095:2026587] = c_w_1343;assign b_s[2028095:2026587] = s_w_1343;
assign b_c[2029604:2028096] = c_w_1344;assign b_s[2029604:2028096] = s_w_1344;
assign b_c[2031113:2029605] = c_w_1345;assign b_s[2031113:2029605] = s_w_1345;
assign b_c[2032622:2031114] = c_w_1346;assign b_s[2032622:2031114] = s_w_1346;
assign b_c[2034131:2032623] = c_w_1347;assign b_s[2034131:2032623] = s_w_1347;
assign b_c[2035640:2034132] = c_w_1348;assign b_s[2035640:2034132] = s_w_1348;
assign b_c[2037149:2035641] = c_w_1349;assign b_s[2037149:2035641] = s_w_1349;
assign b_c[2038658:2037150] = c_w_1350;assign b_s[2038658:2037150] = s_w_1350;
assign b_c[2040167:2038659] = c_w_1351;assign b_s[2040167:2038659] = s_w_1351;
assign b_c[2041676:2040168] = c_w_1352;assign b_s[2041676:2040168] = s_w_1352;
assign b_c[2043185:2041677] = c_w_1353;assign b_s[2043185:2041677] = s_w_1353;
assign b_c[2044694:2043186] = c_w_1354;assign b_s[2044694:2043186] = s_w_1354;
assign b_c[2046203:2044695] = c_w_1355;assign b_s[2046203:2044695] = s_w_1355;
assign b_c[2047712:2046204] = c_w_1356;assign b_s[2047712:2046204] = s_w_1356;
assign b_c[2049221:2047713] = c_w_1357;assign b_s[2049221:2047713] = s_w_1357;
assign b_c[2050730:2049222] = c_w_1358;assign b_s[2050730:2049222] = s_w_1358;
assign b_c[2052239:2050731] = c_w_1359;assign b_s[2052239:2050731] = s_w_1359;
assign b_c[2053748:2052240] = c_w_1360;assign b_s[2053748:2052240] = s_w_1360;
assign b_c[2055257:2053749] = c_w_1361;assign b_s[2055257:2053749] = s_w_1361;
assign b_c[2056766:2055258] = c_w_1362;assign b_s[2056766:2055258] = s_w_1362;
assign b_c[2058275:2056767] = c_w_1363;assign b_s[2058275:2056767] = s_w_1363;
assign b_c[2059784:2058276] = c_w_1364;assign b_s[2059784:2058276] = s_w_1364;
assign b_c[2061293:2059785] = c_w_1365;assign b_s[2061293:2059785] = s_w_1365;
assign b_c[2062802:2061294] = c_w_1366;assign b_s[2062802:2061294] = s_w_1366;
assign b_c[2064311:2062803] = c_w_1367;assign b_s[2064311:2062803] = s_w_1367;
assign b_c[2065820:2064312] = c_w_1368;assign b_s[2065820:2064312] = s_w_1368;
assign b_c[2067329:2065821] = c_w_1369;assign b_s[2067329:2065821] = s_w_1369;
assign b_c[2068838:2067330] = c_w_1370;assign b_s[2068838:2067330] = s_w_1370;
assign b_c[2070347:2068839] = c_w_1371;assign b_s[2070347:2068839] = s_w_1371;
assign b_c[2071856:2070348] = c_w_1372;assign b_s[2071856:2070348] = s_w_1372;
assign b_c[2073365:2071857] = c_w_1373;assign b_s[2073365:2071857] = s_w_1373;
assign b_c[2074874:2073366] = c_w_1374;assign b_s[2074874:2073366] = s_w_1374;
assign b_c[2076383:2074875] = c_w_1375;assign b_s[2076383:2074875] = s_w_1375;
assign b_c[2077892:2076384] = c_w_1376;assign b_s[2077892:2076384] = s_w_1376;
assign b_c[2079401:2077893] = c_w_1377;assign b_s[2079401:2077893] = s_w_1377;
assign b_c[2080910:2079402] = c_w_1378;assign b_s[2080910:2079402] = s_w_1378;
assign b_c[2082419:2080911] = c_w_1379;assign b_s[2082419:2080911] = s_w_1379;
assign b_c[2083928:2082420] = c_w_1380;assign b_s[2083928:2082420] = s_w_1380;
assign b_c[2085437:2083929] = c_w_1381;assign b_s[2085437:2083929] = s_w_1381;
assign b_c[2086946:2085438] = c_w_1382;assign b_s[2086946:2085438] = s_w_1382;
assign b_c[2088455:2086947] = c_w_1383;assign b_s[2088455:2086947] = s_w_1383;
assign b_c[2089964:2088456] = c_w_1384;assign b_s[2089964:2088456] = s_w_1384;
assign b_c[2091473:2089965] = c_w_1385;assign b_s[2091473:2089965] = s_w_1385;
assign b_c[2092982:2091474] = c_w_1386;assign b_s[2092982:2091474] = s_w_1386;
assign b_c[2094491:2092983] = c_w_1387;assign b_s[2094491:2092983] = s_w_1387;
assign b_c[2096000:2094492] = c_w_1388;assign b_s[2096000:2094492] = s_w_1388;
assign b_c[2097509:2096001] = c_w_1389;assign b_s[2097509:2096001] = s_w_1389;
assign b_c[2099018:2097510] = c_w_1390;assign b_s[2099018:2097510] = s_w_1390;
assign b_c[2100527:2099019] = c_w_1391;assign b_s[2100527:2099019] = s_w_1391;
assign b_c[2102036:2100528] = c_w_1392;assign b_s[2102036:2100528] = s_w_1392;
assign b_c[2103545:2102037] = c_w_1393;assign b_s[2103545:2102037] = s_w_1393;
assign b_c[2105054:2103546] = c_w_1394;assign b_s[2105054:2103546] = s_w_1394;
assign b_c[2106563:2105055] = c_w_1395;assign b_s[2106563:2105055] = s_w_1395;
assign b_c[2108072:2106564] = c_w_1396;assign b_s[2108072:2106564] = s_w_1396;
assign b_c[2109581:2108073] = c_w_1397;assign b_s[2109581:2108073] = s_w_1397;
assign b_c[2111090:2109582] = c_w_1398;assign b_s[2111090:2109582] = s_w_1398;
assign b_c[2112599:2111091] = c_w_1399;assign b_s[2112599:2111091] = s_w_1399;
assign b_c[2114108:2112600] = c_w_1400;assign b_s[2114108:2112600] = s_w_1400;
assign b_c[2115617:2114109] = c_w_1401;assign b_s[2115617:2114109] = s_w_1401;
assign b_c[2117126:2115618] = c_w_1402;assign b_s[2117126:2115618] = s_w_1402;
assign b_c[2118635:2117127] = c_w_1403;assign b_s[2118635:2117127] = s_w_1403;
assign b_c[2120144:2118636] = c_w_1404;assign b_s[2120144:2118636] = s_w_1404;
assign b_c[2121653:2120145] = c_w_1405;assign b_s[2121653:2120145] = s_w_1405;
assign b_c[2123162:2121654] = c_w_1406;assign b_s[2123162:2121654] = s_w_1406;
assign b_c[2124671:2123163] = c_w_1407;assign b_s[2124671:2123163] = s_w_1407;
assign b_c[2126180:2124672] = c_w_1408;assign b_s[2126180:2124672] = s_w_1408;
assign b_c[2127689:2126181] = c_w_1409;assign b_s[2127689:2126181] = s_w_1409;
assign b_c[2129198:2127690] = c_w_1410;assign b_s[2129198:2127690] = s_w_1410;
assign b_c[2130707:2129199] = c_w_1411;assign b_s[2130707:2129199] = s_w_1411;
assign b_c[2132216:2130708] = c_w_1412;assign b_s[2132216:2130708] = s_w_1412;
assign b_c[2133725:2132217] = c_w_1413;assign b_s[2133725:2132217] = s_w_1413;
assign b_c[2135234:2133726] = c_w_1414;assign b_s[2135234:2133726] = s_w_1414;
assign b_c[2136743:2135235] = c_w_1415;assign b_s[2136743:2135235] = s_w_1415;
assign b_c[2138252:2136744] = c_w_1416;assign b_s[2138252:2136744] = s_w_1416;
assign b_c[2139761:2138253] = c_w_1417;assign b_s[2139761:2138253] = s_w_1417;
assign b_c[2141270:2139762] = c_w_1418;assign b_s[2141270:2139762] = s_w_1418;
assign b_c[2142779:2141271] = c_w_1419;assign b_s[2142779:2141271] = s_w_1419;
assign b_c[2144288:2142780] = c_w_1420;assign b_s[2144288:2142780] = s_w_1420;
assign b_c[2145797:2144289] = c_w_1421;assign b_s[2145797:2144289] = s_w_1421;
assign b_c[2147306:2145798] = c_w_1422;assign b_s[2147306:2145798] = s_w_1422;
assign b_c[2148815:2147307] = c_w_1423;assign b_s[2148815:2147307] = s_w_1423;
assign b_c[2150324:2148816] = c_w_1424;assign b_s[2150324:2148816] = s_w_1424;
assign b_c[2151833:2150325] = c_w_1425;assign b_s[2151833:2150325] = s_w_1425;
assign b_c[2153342:2151834] = c_w_1426;assign b_s[2153342:2151834] = s_w_1426;
assign b_c[2154851:2153343] = c_w_1427;assign b_s[2154851:2153343] = s_w_1427;
assign b_c[2156360:2154852] = c_w_1428;assign b_s[2156360:2154852] = s_w_1428;
assign b_c[2157869:2156361] = c_w_1429;assign b_s[2157869:2156361] = s_w_1429;
assign b_c[2159378:2157870] = c_w_1430;assign b_s[2159378:2157870] = s_w_1430;
assign b_c[2160887:2159379] = c_w_1431;assign b_s[2160887:2159379] = s_w_1431;
assign b_c[2162396:2160888] = c_w_1432;assign b_s[2162396:2160888] = s_w_1432;
assign b_c[2163905:2162397] = c_w_1433;assign b_s[2163905:2162397] = s_w_1433;
assign b_c[2165414:2163906] = c_w_1434;assign b_s[2165414:2163906] = s_w_1434;
assign b_c[2166923:2165415] = c_w_1435;assign b_s[2166923:2165415] = s_w_1435;
assign b_c[2168432:2166924] = c_w_1436;assign b_s[2168432:2166924] = s_w_1436;
assign b_c[2169941:2168433] = c_w_1437;assign b_s[2169941:2168433] = s_w_1437;
assign b_c[2171450:2169942] = c_w_1438;assign b_s[2171450:2169942] = s_w_1438;
assign b_c[2172959:2171451] = c_w_1439;assign b_s[2172959:2171451] = s_w_1439;
assign b_c[2174468:2172960] = c_w_1440;assign b_s[2174468:2172960] = s_w_1440;
assign b_c[2175977:2174469] = c_w_1441;assign b_s[2175977:2174469] = s_w_1441;
assign b_c[2177486:2175978] = c_w_1442;assign b_s[2177486:2175978] = s_w_1442;
assign b_c[2178995:2177487] = c_w_1443;assign b_s[2178995:2177487] = s_w_1443;
assign b_c[2180504:2178996] = c_w_1444;assign b_s[2180504:2178996] = s_w_1444;
assign b_c[2182013:2180505] = c_w_1445;assign b_s[2182013:2180505] = s_w_1445;
assign b_c[2183522:2182014] = c_w_1446;assign b_s[2183522:2182014] = s_w_1446;
assign b_c[2185031:2183523] = c_w_1447;assign b_s[2185031:2183523] = s_w_1447;
assign b_c[2186540:2185032] = c_w_1448;assign b_s[2186540:2185032] = s_w_1448;
assign b_c[2188049:2186541] = c_w_1449;assign b_s[2188049:2186541] = s_w_1449;
assign b_c[2189558:2188050] = c_w_1450;assign b_s[2189558:2188050] = s_w_1450;
assign b_c[2191067:2189559] = c_w_1451;assign b_s[2191067:2189559] = s_w_1451;
assign b_c[2192576:2191068] = c_w_1452;assign b_s[2192576:2191068] = s_w_1452;
assign b_c[2194085:2192577] = c_w_1453;assign b_s[2194085:2192577] = s_w_1453;
assign b_c[2195594:2194086] = c_w_1454;assign b_s[2195594:2194086] = s_w_1454;
assign b_c[2197103:2195595] = c_w_1455;assign b_s[2197103:2195595] = s_w_1455;
assign b_c[2198612:2197104] = c_w_1456;assign b_s[2198612:2197104] = s_w_1456;
assign b_c[2200121:2198613] = c_w_1457;assign b_s[2200121:2198613] = s_w_1457;
assign b_c[2201630:2200122] = c_w_1458;assign b_s[2201630:2200122] = s_w_1458;
assign b_c[2203139:2201631] = c_w_1459;assign b_s[2203139:2201631] = s_w_1459;
assign b_c[2204648:2203140] = c_w_1460;assign b_s[2204648:2203140] = s_w_1460;
assign b_c[2206157:2204649] = c_w_1461;assign b_s[2206157:2204649] = s_w_1461;
assign b_c[2207666:2206158] = c_w_1462;assign b_s[2207666:2206158] = s_w_1462;
assign b_c[2209175:2207667] = c_w_1463;assign b_s[2209175:2207667] = s_w_1463;
assign b_c[2210684:2209176] = c_w_1464;assign b_s[2210684:2209176] = s_w_1464;
assign b_c[2212193:2210685] = c_w_1465;assign b_s[2212193:2210685] = s_w_1465;
assign b_c[2213702:2212194] = c_w_1466;assign b_s[2213702:2212194] = s_w_1466;
assign b_c[2215211:2213703] = c_w_1467;assign b_s[2215211:2213703] = s_w_1467;
assign b_c[2216720:2215212] = c_w_1468;assign b_s[2216720:2215212] = s_w_1468;
assign b_c[2218229:2216721] = c_w_1469;assign b_s[2218229:2216721] = s_w_1469;
assign b_c[2219738:2218230] = c_w_1470;assign b_s[2219738:2218230] = s_w_1470;
assign b_c[2221247:2219739] = c_w_1471;assign b_s[2221247:2219739] = s_w_1471;
assign b_c[2222756:2221248] = c_w_1472;assign b_s[2222756:2221248] = s_w_1472;
assign b_c[2224265:2222757] = c_w_1473;assign b_s[2224265:2222757] = s_w_1473;
assign b_c[2225774:2224266] = c_w_1474;assign b_s[2225774:2224266] = s_w_1474;
assign b_c[2227283:2225775] = c_w_1475;assign b_s[2227283:2225775] = s_w_1475;
assign b_c[2228792:2227284] = c_w_1476;assign b_s[2228792:2227284] = s_w_1476;
assign b_c[2230301:2228793] = c_w_1477;assign b_s[2230301:2228793] = s_w_1477;
assign b_c[2231810:2230302] = c_w_1478;assign b_s[2231810:2230302] = s_w_1478;
assign b_c[2233319:2231811] = c_w_1479;assign b_s[2233319:2231811] = s_w_1479;
assign b_c[2234828:2233320] = c_w_1480;assign b_s[2234828:2233320] = s_w_1480;
assign b_c[2236337:2234829] = c_w_1481;assign b_s[2236337:2234829] = s_w_1481;
assign b_c[2237846:2236338] = c_w_1482;assign b_s[2237846:2236338] = s_w_1482;
assign b_c[2239355:2237847] = c_w_1483;assign b_s[2239355:2237847] = s_w_1483;
assign b_c[2240864:2239356] = c_w_1484;assign b_s[2240864:2239356] = s_w_1484;
assign b_c[2242373:2240865] = c_w_1485;assign b_s[2242373:2240865] = s_w_1485;
assign b_c[2243882:2242374] = c_w_1486;assign b_s[2243882:2242374] = s_w_1486;
assign b_c[2245391:2243883] = c_w_1487;assign b_s[2245391:2243883] = s_w_1487;
assign b_c[2246900:2245392] = c_w_1488;assign b_s[2246900:2245392] = s_w_1488;
assign b_c[2248409:2246901] = c_w_1489;assign b_s[2248409:2246901] = s_w_1489;
assign b_c[2249918:2248410] = c_w_1490;assign b_s[2249918:2248410] = s_w_1490;
assign b_c[2251427:2249919] = c_w_1491;assign b_s[2251427:2249919] = s_w_1491;
assign b_c[2252936:2251428] = c_w_1492;assign b_s[2252936:2251428] = s_w_1492;
assign b_c[2254445:2252937] = c_w_1493;assign b_s[2254445:2252937] = s_w_1493;
assign b_c[2255954:2254446] = c_w_1494;assign b_s[2255954:2254446] = s_w_1494;
assign b_c[2257463:2255955] = c_w_1495;assign b_s[2257463:2255955] = s_w_1495;
assign b_c[2258972:2257464] = c_w_1496;assign b_s[2258972:2257464] = s_w_1496;
assign b_c[2260481:2258973] = c_w_1497;assign b_s[2260481:2258973] = s_w_1497;
assign b_c[2261990:2260482] = c_w_1498;assign b_s[2261990:2260482] = s_w_1498;
assign b_c[2263499:2261991] = c_w_1499;assign b_s[2263499:2261991] = s_w_1499;
assign b_c[2265008:2263500] = c_w_1500;assign b_s[2265008:2263500] = s_w_1500;
assign b_c[2266517:2265009] = c_w_1501;assign b_s[2266517:2265009] = s_w_1501;
assign b_c[2268026:2266518] = c_w_1502;assign b_s[2268026:2266518] = s_w_1502;
assign b_c[2269535:2268027] = c_w_1503;assign b_s[2269535:2268027] = s_w_1503;
assign b_c[2271044:2269536] = c_w_1504;assign b_s[2271044:2269536] = s_w_1504;
assign b_c[2272553:2271045] = c_w_1505;assign b_s[2272553:2271045] = s_w_1505;
assign b_c[2274062:2272554] = c_w_1506;assign b_s[2274062:2272554] = s_w_1506;
assign b_c[2275571:2274063] = c_w_1507;assign b_s[2275571:2274063] = s_w_1507;
assign b_c[2277080:2275572] = c_w_1508;assign b_s[2277080:2275572] = s_w_1508;
    
endmodule
    