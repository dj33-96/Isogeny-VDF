
module xor_40_array(
    input [39:0] in0,in1,
    output [39:0] out0
);

assign out0 = in0 ^ in1;

endmodule
    