

module csa_tree_89x178(
    input [15841:0] A, // lines are appended together
    output[177:0] B_0,
    output[177:0] B_1
);

wire [10679:0] tree_1;
wire [7119:0] tree_2;
wire [4805:0] tree_3;
wire [3203:0] tree_4;
wire [2135:0] tree_5;
wire [1423:0] tree_6;
wire [1067:0] tree_7;
wire [711:0] tree_8;
wire [533:0] tree_9;
wire [355:0] tree_10;
// layer-1
csa_178 csau_178_i0(A[177:0],A[355:178],A[533:356],tree_1[177:0],tree_1[355:178]);
csa_178 csau_178_i1(A[711:534],A[889:712],A[1067:890],tree_1[533:356],tree_1[711:534]);
csa_178 csau_178_i2(A[1245:1068],A[1423:1246],A[1601:1424],tree_1[889:712],tree_1[1067:890]);
csa_178 csau_178_i3(A[1779:1602],A[1957:1780],A[2135:1958],tree_1[1245:1068],tree_1[1423:1246]);
csa_178 csau_178_i4(A[2313:2136],A[2491:2314],A[2669:2492],tree_1[1601:1424],tree_1[1779:1602]);
csa_178 csau_178_i5(A[2847:2670],A[3025:2848],A[3203:3026],tree_1[1957:1780],tree_1[2135:1958]);
csa_178 csau_178_i6(A[3381:3204],A[3559:3382],A[3737:3560],tree_1[2313:2136],tree_1[2491:2314]);
csa_178 csau_178_i7(A[3915:3738],A[4093:3916],A[4271:4094],tree_1[2669:2492],tree_1[2847:2670]);
csa_178 csau_178_i8(A[4449:4272],A[4627:4450],A[4805:4628],tree_1[3025:2848],tree_1[3203:3026]);
csa_178 csau_178_i9(A[4983:4806],A[5161:4984],A[5339:5162],tree_1[3381:3204],tree_1[3559:3382]);
csa_178 csau_178_i10(A[5517:5340],A[5695:5518],A[5873:5696],tree_1[3737:3560],tree_1[3915:3738]);
csa_178 csau_178_i11(A[6051:5874],A[6229:6052],A[6407:6230],tree_1[4093:3916],tree_1[4271:4094]);
csa_178 csau_178_i12(A[6585:6408],A[6763:6586],A[6941:6764],tree_1[4449:4272],tree_1[4627:4450]);
csa_178 csau_178_i13(A[7119:6942],A[7297:7120],A[7475:7298],tree_1[4805:4628],tree_1[4983:4806]);
csa_178 csau_178_i14(A[7653:7476],A[7831:7654],A[8009:7832],tree_1[5161:4984],tree_1[5339:5162]);
csa_178 csau_178_i15(A[8187:8010],A[8365:8188],A[8543:8366],tree_1[5517:5340],tree_1[5695:5518]);
csa_178 csau_178_i16(A[8721:8544],A[8899:8722],A[9077:8900],tree_1[5873:5696],tree_1[6051:5874]);
csa_178 csau_178_i17(A[9255:9078],A[9433:9256],A[9611:9434],tree_1[6229:6052],tree_1[6407:6230]);
csa_178 csau_178_i18(A[9789:9612],A[9967:9790],A[10145:9968],tree_1[6585:6408],tree_1[6763:6586]);
csa_178 csau_178_i19(A[10323:10146],A[10501:10324],A[10679:10502],tree_1[6941:6764],tree_1[7119:6942]);
csa_178 csau_178_i20(A[10857:10680],A[11035:10858],A[11213:11036],tree_1[7297:7120],tree_1[7475:7298]);
csa_178 csau_178_i21(A[11391:11214],A[11569:11392],A[11747:11570],tree_1[7653:7476],tree_1[7831:7654]);
csa_178 csau_178_i22(A[11925:11748],A[12103:11926],A[12281:12104],tree_1[8009:7832],tree_1[8187:8010]);
csa_178 csau_178_i23(A[12459:12282],A[12637:12460],A[12815:12638],tree_1[8365:8188],tree_1[8543:8366]);
csa_178 csau_178_i24(A[12993:12816],A[13171:12994],A[13349:13172],tree_1[8721:8544],tree_1[8899:8722]);
csa_178 csau_178_i25(A[13527:13350],A[13705:13528],A[13883:13706],tree_1[9077:8900],tree_1[9255:9078]);
csa_178 csau_178_i26(A[14061:13884],A[14239:14062],A[14417:14240],tree_1[9433:9256],tree_1[9611:9434]);
csa_178 csau_178_i27(A[14595:14418],A[14773:14596],A[14951:14774],tree_1[9789:9612],tree_1[9967:9790]);
csa_178 csau_178_i28(A[15129:14952],A[15307:15130],A[15485:15308],tree_1[10145:9968],tree_1[10323:10146]);
assign tree_1[10501:10324] = A[15663:15486];
assign tree_1[10679:10502] = A[15841:15664];
// layer-2
csa_178 csau_178_i29(tree_1[177:0],tree_1[355:178],tree_1[533:356],tree_2[177:0],tree_2[355:178]);
csa_178 csau_178_i30(tree_1[711:534],tree_1[889:712],tree_1[1067:890],tree_2[533:356],tree_2[711:534]);
csa_178 csau_178_i31(tree_1[1245:1068],tree_1[1423:1246],tree_1[1601:1424],tree_2[889:712],tree_2[1067:890]);
csa_178 csau_178_i32(tree_1[1779:1602],tree_1[1957:1780],tree_1[2135:1958],tree_2[1245:1068],tree_2[1423:1246]);
csa_178 csau_178_i33(tree_1[2313:2136],tree_1[2491:2314],tree_1[2669:2492],tree_2[1601:1424],tree_2[1779:1602]);
csa_178 csau_178_i34(tree_1[2847:2670],tree_1[3025:2848],tree_1[3203:3026],tree_2[1957:1780],tree_2[2135:1958]);
csa_178 csau_178_i35(tree_1[3381:3204],tree_1[3559:3382],tree_1[3737:3560],tree_2[2313:2136],tree_2[2491:2314]);
csa_178 csau_178_i36(tree_1[3915:3738],tree_1[4093:3916],tree_1[4271:4094],tree_2[2669:2492],tree_2[2847:2670]);
csa_178 csau_178_i37(tree_1[4449:4272],tree_1[4627:4450],tree_1[4805:4628],tree_2[3025:2848],tree_2[3203:3026]);
csa_178 csau_178_i38(tree_1[4983:4806],tree_1[5161:4984],tree_1[5339:5162],tree_2[3381:3204],tree_2[3559:3382]);
csa_178 csau_178_i39(tree_1[5517:5340],tree_1[5695:5518],tree_1[5873:5696],tree_2[3737:3560],tree_2[3915:3738]);
csa_178 csau_178_i40(tree_1[6051:5874],tree_1[6229:6052],tree_1[6407:6230],tree_2[4093:3916],tree_2[4271:4094]);
csa_178 csau_178_i41(tree_1[6585:6408],tree_1[6763:6586],tree_1[6941:6764],tree_2[4449:4272],tree_2[4627:4450]);
csa_178 csau_178_i42(tree_1[7119:6942],tree_1[7297:7120],tree_1[7475:7298],tree_2[4805:4628],tree_2[4983:4806]);
csa_178 csau_178_i43(tree_1[7653:7476],tree_1[7831:7654],tree_1[8009:7832],tree_2[5161:4984],tree_2[5339:5162]);
csa_178 csau_178_i44(tree_1[8187:8010],tree_1[8365:8188],tree_1[8543:8366],tree_2[5517:5340],tree_2[5695:5518]);
csa_178 csau_178_i45(tree_1[8721:8544],tree_1[8899:8722],tree_1[9077:8900],tree_2[5873:5696],tree_2[6051:5874]);
csa_178 csau_178_i46(tree_1[9255:9078],tree_1[9433:9256],tree_1[9611:9434],tree_2[6229:6052],tree_2[6407:6230]);
csa_178 csau_178_i47(tree_1[9789:9612],tree_1[9967:9790],tree_1[10145:9968],tree_2[6585:6408],tree_2[6763:6586]);
csa_178 csau_178_i48(tree_1[10323:10146],tree_1[10501:10324],tree_1[10679:10502],tree_2[6941:6764],tree_2[7119:6942]);
// layer-3
csa_178 csau_178_i49(tree_2[177:0],tree_2[355:178],tree_2[533:356],tree_3[177:0],tree_3[355:178]);
csa_178 csau_178_i50(tree_2[711:534],tree_2[889:712],tree_2[1067:890],tree_3[533:356],tree_3[711:534]);
csa_178 csau_178_i51(tree_2[1245:1068],tree_2[1423:1246],tree_2[1601:1424],tree_3[889:712],tree_3[1067:890]);
csa_178 csau_178_i52(tree_2[1779:1602],tree_2[1957:1780],tree_2[2135:1958],tree_3[1245:1068],tree_3[1423:1246]);
csa_178 csau_178_i53(tree_2[2313:2136],tree_2[2491:2314],tree_2[2669:2492],tree_3[1601:1424],tree_3[1779:1602]);
csa_178 csau_178_i54(tree_2[2847:2670],tree_2[3025:2848],tree_2[3203:3026],tree_3[1957:1780],tree_3[2135:1958]);
csa_178 csau_178_i55(tree_2[3381:3204],tree_2[3559:3382],tree_2[3737:3560],tree_3[2313:2136],tree_3[2491:2314]);
csa_178 csau_178_i56(tree_2[3915:3738],tree_2[4093:3916],tree_2[4271:4094],tree_3[2669:2492],tree_3[2847:2670]);
csa_178 csau_178_i57(tree_2[4449:4272],tree_2[4627:4450],tree_2[4805:4628],tree_3[3025:2848],tree_3[3203:3026]);
csa_178 csau_178_i58(tree_2[4983:4806],tree_2[5161:4984],tree_2[5339:5162],tree_3[3381:3204],tree_3[3559:3382]);
csa_178 csau_178_i59(tree_2[5517:5340],tree_2[5695:5518],tree_2[5873:5696],tree_3[3737:3560],tree_3[3915:3738]);
csa_178 csau_178_i60(tree_2[6051:5874],tree_2[6229:6052],tree_2[6407:6230],tree_3[4093:3916],tree_3[4271:4094]);
csa_178 csau_178_i61(tree_2[6585:6408],tree_2[6763:6586],tree_2[6941:6764],tree_3[4449:4272],tree_3[4627:4450]);
assign tree_3[4805:4628] = tree_2[7119:6942];
// layer-4
csa_178 csau_178_i62(tree_3[177:0],tree_3[355:178],tree_3[533:356],tree_4[177:0],tree_4[355:178]);
csa_178 csau_178_i63(tree_3[711:534],tree_3[889:712],tree_3[1067:890],tree_4[533:356],tree_4[711:534]);
csa_178 csau_178_i64(tree_3[1245:1068],tree_3[1423:1246],tree_3[1601:1424],tree_4[889:712],tree_4[1067:890]);
csa_178 csau_178_i65(tree_3[1779:1602],tree_3[1957:1780],tree_3[2135:1958],tree_4[1245:1068],tree_4[1423:1246]);
csa_178 csau_178_i66(tree_3[2313:2136],tree_3[2491:2314],tree_3[2669:2492],tree_4[1601:1424],tree_4[1779:1602]);
csa_178 csau_178_i67(tree_3[2847:2670],tree_3[3025:2848],tree_3[3203:3026],tree_4[1957:1780],tree_4[2135:1958]);
csa_178 csau_178_i68(tree_3[3381:3204],tree_3[3559:3382],tree_3[3737:3560],tree_4[2313:2136],tree_4[2491:2314]);
csa_178 csau_178_i69(tree_3[3915:3738],tree_3[4093:3916],tree_3[4271:4094],tree_4[2669:2492],tree_4[2847:2670]);
csa_178 csau_178_i70(tree_3[4449:4272],tree_3[4627:4450],tree_3[4805:4628],tree_4[3025:2848],tree_4[3203:3026]);
// layer-5
csa_178 csau_178_i71(tree_4[177:0],tree_4[355:178],tree_4[533:356],tree_5[177:0],tree_5[355:178]);
csa_178 csau_178_i72(tree_4[711:534],tree_4[889:712],tree_4[1067:890],tree_5[533:356],tree_5[711:534]);
csa_178 csau_178_i73(tree_4[1245:1068],tree_4[1423:1246],tree_4[1601:1424],tree_5[889:712],tree_5[1067:890]);
csa_178 csau_178_i74(tree_4[1779:1602],tree_4[1957:1780],tree_4[2135:1958],tree_5[1245:1068],tree_5[1423:1246]);
csa_178 csau_178_i75(tree_4[2313:2136],tree_4[2491:2314],tree_4[2669:2492],tree_5[1601:1424],tree_5[1779:1602]);
csa_178 csau_178_i76(tree_4[2847:2670],tree_4[3025:2848],tree_4[3203:3026],tree_5[1957:1780],tree_5[2135:1958]);
// layer-6
csa_178 csau_178_i77(tree_5[177:0],tree_5[355:178],tree_5[533:356],tree_6[177:0],tree_6[355:178]);
csa_178 csau_178_i78(tree_5[711:534],tree_5[889:712],tree_5[1067:890],tree_6[533:356],tree_6[711:534]);
csa_178 csau_178_i79(tree_5[1245:1068],tree_5[1423:1246],tree_5[1601:1424],tree_6[889:712],tree_6[1067:890]);
csa_178 csau_178_i80(tree_5[1779:1602],tree_5[1957:1780],tree_5[2135:1958],tree_6[1245:1068],tree_6[1423:1246]);
// layer-7
csa_178 csau_178_i81(tree_6[177:0],tree_6[355:178],tree_6[533:356],tree_7[177:0],tree_7[355:178]);
csa_178 csau_178_i82(tree_6[711:534],tree_6[889:712],tree_6[1067:890],tree_7[533:356],tree_7[711:534]);
assign tree_7[889:712] = tree_6[1245:1068];
assign tree_7[1067:890] = tree_6[1423:1246];
// layer-8
csa_178 csau_178_i83(tree_7[177:0],tree_7[355:178],tree_7[533:356],tree_8[177:0],tree_8[355:178]);
csa_178 csau_178_i84(tree_7[711:534],tree_7[889:712],tree_7[1067:890],tree_8[533:356],tree_8[711:534]);
// layer-9
csa_178 csau_178_i85(tree_8[177:0],tree_8[355:178],tree_8[533:356],tree_9[177:0],tree_9[355:178]);
assign tree_9[533:356] = tree_8[711:534];
// layer-10
csa_178 csau_178_i86(tree_9[177:0],tree_9[355:178],tree_9[533:356],tree_10[177:0],tree_10[355:178]);

// final assignment
assign B_0 = tree_10[177:0];
assign B_1 = tree_10[355:178];

endmodule
