
module csa_80 (
    input [79:0] x,y,z,
    output[79:0] c,s 
);

wire dummy;

assign c[0] = 1'b0;
    
assign {c[1],s[0]} = (x[0]+y[0]+z[0]);
assign {c[2],s[1]} = (x[1]+y[1]+z[1]);
assign {c[3],s[2]} = (x[2]+y[2]+z[2]);
assign {c[4],s[3]} = (x[3]+y[3]+z[3]);
assign {c[5],s[4]} = (x[4]+y[4]+z[4]);
assign {c[6],s[5]} = (x[5]+y[5]+z[5]);
assign {c[7],s[6]} = (x[6]+y[6]+z[6]);
assign {c[8],s[7]} = (x[7]+y[7]+z[7]);
assign {c[9],s[8]} = (x[8]+y[8]+z[8]);
assign {c[10],s[9]} = (x[9]+y[9]+z[9]);
assign {c[11],s[10]} = (x[10]+y[10]+z[10]);
assign {c[12],s[11]} = (x[11]+y[11]+z[11]);
assign {c[13],s[12]} = (x[12]+y[12]+z[12]);
assign {c[14],s[13]} = (x[13]+y[13]+z[13]);
assign {c[15],s[14]} = (x[14]+y[14]+z[14]);
assign {c[16],s[15]} = (x[15]+y[15]+z[15]);
assign {c[17],s[16]} = (x[16]+y[16]+z[16]);
assign {c[18],s[17]} = (x[17]+y[17]+z[17]);
assign {c[19],s[18]} = (x[18]+y[18]+z[18]);
assign {c[20],s[19]} = (x[19]+y[19]+z[19]);
assign {c[21],s[20]} = (x[20]+y[20]+z[20]);
assign {c[22],s[21]} = (x[21]+y[21]+z[21]);
assign {c[23],s[22]} = (x[22]+y[22]+z[22]);
assign {c[24],s[23]} = (x[23]+y[23]+z[23]);
assign {c[25],s[24]} = (x[24]+y[24]+z[24]);
assign {c[26],s[25]} = (x[25]+y[25]+z[25]);
assign {c[27],s[26]} = (x[26]+y[26]+z[26]);
assign {c[28],s[27]} = (x[27]+y[27]+z[27]);
assign {c[29],s[28]} = (x[28]+y[28]+z[28]);
assign {c[30],s[29]} = (x[29]+y[29]+z[29]);
assign {c[31],s[30]} = (x[30]+y[30]+z[30]);
assign {c[32],s[31]} = (x[31]+y[31]+z[31]);
assign {c[33],s[32]} = (x[32]+y[32]+z[32]);
assign {c[34],s[33]} = (x[33]+y[33]+z[33]);
assign {c[35],s[34]} = (x[34]+y[34]+z[34]);
assign {c[36],s[35]} = (x[35]+y[35]+z[35]);
assign {c[37],s[36]} = (x[36]+y[36]+z[36]);
assign {c[38],s[37]} = (x[37]+y[37]+z[37]);
assign {c[39],s[38]} = (x[38]+y[38]+z[38]);
assign {c[40],s[39]} = (x[39]+y[39]+z[39]);
assign {c[41],s[40]} = (x[40]+y[40]+z[40]);
assign {c[42],s[41]} = (x[41]+y[41]+z[41]);
assign {c[43],s[42]} = (x[42]+y[42]+z[42]);
assign {c[44],s[43]} = (x[43]+y[43]+z[43]);
assign {c[45],s[44]} = (x[44]+y[44]+z[44]);
assign {c[46],s[45]} = (x[45]+y[45]+z[45]);
assign {c[47],s[46]} = (x[46]+y[46]+z[46]);
assign {c[48],s[47]} = (x[47]+y[47]+z[47]);
assign {c[49],s[48]} = (x[48]+y[48]+z[48]);
assign {c[50],s[49]} = (x[49]+y[49]+z[49]);
assign {c[51],s[50]} = (x[50]+y[50]+z[50]);
assign {c[52],s[51]} = (x[51]+y[51]+z[51]);
assign {c[53],s[52]} = (x[52]+y[52]+z[52]);
assign {c[54],s[53]} = (x[53]+y[53]+z[53]);
assign {c[55],s[54]} = (x[54]+y[54]+z[54]);
assign {c[56],s[55]} = (x[55]+y[55]+z[55]);
assign {c[57],s[56]} = (x[56]+y[56]+z[56]);
assign {c[58],s[57]} = (x[57]+y[57]+z[57]);
assign {c[59],s[58]} = (x[58]+y[58]+z[58]);
assign {c[60],s[59]} = (x[59]+y[59]+z[59]);
assign {c[61],s[60]} = (x[60]+y[60]+z[60]);
assign {c[62],s[61]} = (x[61]+y[61]+z[61]);
assign {c[63],s[62]} = (x[62]+y[62]+z[62]);
assign {c[64],s[63]} = (x[63]+y[63]+z[63]);
assign {c[65],s[64]} = (x[64]+y[64]+z[64]);
assign {c[66],s[65]} = (x[65]+y[65]+z[65]);
assign {c[67],s[66]} = (x[66]+y[66]+z[66]);
assign {c[68],s[67]} = (x[67]+y[67]+z[67]);
assign {c[69],s[68]} = (x[68]+y[68]+z[68]);
assign {c[70],s[69]} = (x[69]+y[69]+z[69]);
assign {c[71],s[70]} = (x[70]+y[70]+z[70]);
assign {c[72],s[71]} = (x[71]+y[71]+z[71]);
assign {c[73],s[72]} = (x[72]+y[72]+z[72]);
assign {c[74],s[73]} = (x[73]+y[73]+z[73]);
assign {c[75],s[74]} = (x[74]+y[74]+z[74]);
assign {c[76],s[75]} = (x[75]+y[75]+z[75]);
assign {c[77],s[76]} = (x[76]+y[76]+z[76]);
assign {c[78],s[77]} = (x[77]+y[77]+z[77]);
assign {c[79],s[78]} = (x[78]+y[78]+z[78]);
assign {dummy,s[79]} = (x[79]+y[79]+z[79]);

endmodule
    