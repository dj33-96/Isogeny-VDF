
module AND_matrix_92x92(
    input [91:0] a,
    input [91:0] b,
    output [16927:0] c // lines are appended together
);
    
wire [91:0] c_w_0;
wire [91:0] c_w_1;
wire [91:0] c_w_2;
wire [91:0] c_w_3;
wire [91:0] c_w_4;
wire [91:0] c_w_5;
wire [91:0] c_w_6;
wire [91:0] c_w_7;
wire [91:0] c_w_8;
wire [91:0] c_w_9;
wire [91:0] c_w_10;
wire [91:0] c_w_11;
wire [91:0] c_w_12;
wire [91:0] c_w_13;
wire [91:0] c_w_14;
wire [91:0] c_w_15;
wire [91:0] c_w_16;
wire [91:0] c_w_17;
wire [91:0] c_w_18;
wire [91:0] c_w_19;
wire [91:0] c_w_20;
wire [91:0] c_w_21;
wire [91:0] c_w_22;
wire [91:0] c_w_23;
wire [91:0] c_w_24;
wire [91:0] c_w_25;
wire [91:0] c_w_26;
wire [91:0] c_w_27;
wire [91:0] c_w_28;
wire [91:0] c_w_29;
wire [91:0] c_w_30;
wire [91:0] c_w_31;
wire [91:0] c_w_32;
wire [91:0] c_w_33;
wire [91:0] c_w_34;
wire [91:0] c_w_35;
wire [91:0] c_w_36;
wire [91:0] c_w_37;
wire [91:0] c_w_38;
wire [91:0] c_w_39;
wire [91:0] c_w_40;
wire [91:0] c_w_41;
wire [91:0] c_w_42;
wire [91:0] c_w_43;
wire [91:0] c_w_44;
wire [91:0] c_w_45;
wire [91:0] c_w_46;
wire [91:0] c_w_47;
wire [91:0] c_w_48;
wire [91:0] c_w_49;
wire [91:0] c_w_50;
wire [91:0] c_w_51;
wire [91:0] c_w_52;
wire [91:0] c_w_53;
wire [91:0] c_w_54;
wire [91:0] c_w_55;
wire [91:0] c_w_56;
wire [91:0] c_w_57;
wire [91:0] c_w_58;
wire [91:0] c_w_59;
wire [91:0] c_w_60;
wire [91:0] c_w_61;
wire [91:0] c_w_62;
wire [91:0] c_w_63;
wire [91:0] c_w_64;
wire [91:0] c_w_65;
wire [91:0] c_w_66;
wire [91:0] c_w_67;
wire [91:0] c_w_68;
wire [91:0] c_w_69;
wire [91:0] c_w_70;
wire [91:0] c_w_71;
wire [91:0] c_w_72;
wire [91:0] c_w_73;
wire [91:0] c_w_74;
wire [91:0] c_w_75;
wire [91:0] c_w_76;
wire [91:0] c_w_77;
wire [91:0] c_w_78;
wire [91:0] c_w_79;
wire [91:0] c_w_80;
wire [91:0] c_w_81;
wire [91:0] c_w_82;
wire [91:0] c_w_83;
wire [91:0] c_w_84;
wire [91:0] c_w_85;
wire [91:0] c_w_86;
wire [91:0] c_w_87;
wire [91:0] c_w_88;
wire [91:0] c_w_89;
wire [91:0] c_w_90;
wire [91:0] c_w_91;
    
AND_array_92 AND_array_92_i0(a,b[0],c_w_0);
AND_array_92 AND_array_92_i1(a,b[1],c_w_1);
AND_array_92 AND_array_92_i2(a,b[2],c_w_2);
AND_array_92 AND_array_92_i3(a,b[3],c_w_3);
AND_array_92 AND_array_92_i4(a,b[4],c_w_4);
AND_array_92 AND_array_92_i5(a,b[5],c_w_5);
AND_array_92 AND_array_92_i6(a,b[6],c_w_6);
AND_array_92 AND_array_92_i7(a,b[7],c_w_7);
AND_array_92 AND_array_92_i8(a,b[8],c_w_8);
AND_array_92 AND_array_92_i9(a,b[9],c_w_9);
AND_array_92 AND_array_92_i10(a,b[10],c_w_10);
AND_array_92 AND_array_92_i11(a,b[11],c_w_11);
AND_array_92 AND_array_92_i12(a,b[12],c_w_12);
AND_array_92 AND_array_92_i13(a,b[13],c_w_13);
AND_array_92 AND_array_92_i14(a,b[14],c_w_14);
AND_array_92 AND_array_92_i15(a,b[15],c_w_15);
AND_array_92 AND_array_92_i16(a,b[16],c_w_16);
AND_array_92 AND_array_92_i17(a,b[17],c_w_17);
AND_array_92 AND_array_92_i18(a,b[18],c_w_18);
AND_array_92 AND_array_92_i19(a,b[19],c_w_19);
AND_array_92 AND_array_92_i20(a,b[20],c_w_20);
AND_array_92 AND_array_92_i21(a,b[21],c_w_21);
AND_array_92 AND_array_92_i22(a,b[22],c_w_22);
AND_array_92 AND_array_92_i23(a,b[23],c_w_23);
AND_array_92 AND_array_92_i24(a,b[24],c_w_24);
AND_array_92 AND_array_92_i25(a,b[25],c_w_25);
AND_array_92 AND_array_92_i26(a,b[26],c_w_26);
AND_array_92 AND_array_92_i27(a,b[27],c_w_27);
AND_array_92 AND_array_92_i28(a,b[28],c_w_28);
AND_array_92 AND_array_92_i29(a,b[29],c_w_29);
AND_array_92 AND_array_92_i30(a,b[30],c_w_30);
AND_array_92 AND_array_92_i31(a,b[31],c_w_31);
AND_array_92 AND_array_92_i32(a,b[32],c_w_32);
AND_array_92 AND_array_92_i33(a,b[33],c_w_33);
AND_array_92 AND_array_92_i34(a,b[34],c_w_34);
AND_array_92 AND_array_92_i35(a,b[35],c_w_35);
AND_array_92 AND_array_92_i36(a,b[36],c_w_36);
AND_array_92 AND_array_92_i37(a,b[37],c_w_37);
AND_array_92 AND_array_92_i38(a,b[38],c_w_38);
AND_array_92 AND_array_92_i39(a,b[39],c_w_39);
AND_array_92 AND_array_92_i40(a,b[40],c_w_40);
AND_array_92 AND_array_92_i41(a,b[41],c_w_41);
AND_array_92 AND_array_92_i42(a,b[42],c_w_42);
AND_array_92 AND_array_92_i43(a,b[43],c_w_43);
AND_array_92 AND_array_92_i44(a,b[44],c_w_44);
AND_array_92 AND_array_92_i45(a,b[45],c_w_45);
AND_array_92 AND_array_92_i46(a,b[46],c_w_46);
AND_array_92 AND_array_92_i47(a,b[47],c_w_47);
AND_array_92 AND_array_92_i48(a,b[48],c_w_48);
AND_array_92 AND_array_92_i49(a,b[49],c_w_49);
AND_array_92 AND_array_92_i50(a,b[50],c_w_50);
AND_array_92 AND_array_92_i51(a,b[51],c_w_51);
AND_array_92 AND_array_92_i52(a,b[52],c_w_52);
AND_array_92 AND_array_92_i53(a,b[53],c_w_53);
AND_array_92 AND_array_92_i54(a,b[54],c_w_54);
AND_array_92 AND_array_92_i55(a,b[55],c_w_55);
AND_array_92 AND_array_92_i56(a,b[56],c_w_56);
AND_array_92 AND_array_92_i57(a,b[57],c_w_57);
AND_array_92 AND_array_92_i58(a,b[58],c_w_58);
AND_array_92 AND_array_92_i59(a,b[59],c_w_59);
AND_array_92 AND_array_92_i60(a,b[60],c_w_60);
AND_array_92 AND_array_92_i61(a,b[61],c_w_61);
AND_array_92 AND_array_92_i62(a,b[62],c_w_62);
AND_array_92 AND_array_92_i63(a,b[63],c_w_63);
AND_array_92 AND_array_92_i64(a,b[64],c_w_64);
AND_array_92 AND_array_92_i65(a,b[65],c_w_65);
AND_array_92 AND_array_92_i66(a,b[66],c_w_66);
AND_array_92 AND_array_92_i67(a,b[67],c_w_67);
AND_array_92 AND_array_92_i68(a,b[68],c_w_68);
AND_array_92 AND_array_92_i69(a,b[69],c_w_69);
AND_array_92 AND_array_92_i70(a,b[70],c_w_70);
AND_array_92 AND_array_92_i71(a,b[71],c_w_71);
AND_array_92 AND_array_92_i72(a,b[72],c_w_72);
AND_array_92 AND_array_92_i73(a,b[73],c_w_73);
AND_array_92 AND_array_92_i74(a,b[74],c_w_74);
AND_array_92 AND_array_92_i75(a,b[75],c_w_75);
AND_array_92 AND_array_92_i76(a,b[76],c_w_76);
AND_array_92 AND_array_92_i77(a,b[77],c_w_77);
AND_array_92 AND_array_92_i78(a,b[78],c_w_78);
AND_array_92 AND_array_92_i79(a,b[79],c_w_79);
AND_array_92 AND_array_92_i80(a,b[80],c_w_80);
AND_array_92 AND_array_92_i81(a,b[81],c_w_81);
AND_array_92 AND_array_92_i82(a,b[82],c_w_82);
AND_array_92 AND_array_92_i83(a,b[83],c_w_83);
AND_array_92 AND_array_92_i84(a,b[84],c_w_84);
AND_array_92 AND_array_92_i85(a,b[85],c_w_85);
AND_array_92 AND_array_92_i86(a,b[86],c_w_86);
AND_array_92 AND_array_92_i87(a,b[87],c_w_87);
AND_array_92 AND_array_92_i88(a,b[88],c_w_88);
AND_array_92 AND_array_92_i89(a,b[89],c_w_89);
AND_array_92 AND_array_92_i90(a,b[90],c_w_90);
AND_array_92 AND_array_92_i91(a,b[91],c_w_91);
    
assign c[183:0] = {92'b0,c_w_0};
assign c[367:184] = {91'b0,c_w_1,1'b0};
assign c[551:368] = {90'b0,c_w_2,2'b0};
assign c[735:552] = {89'b0,c_w_3,3'b0};
assign c[919:736] = {88'b0,c_w_4,4'b0};
assign c[1103:920] = {87'b0,c_w_5,5'b0};
assign c[1287:1104] = {86'b0,c_w_6,6'b0};
assign c[1471:1288] = {85'b0,c_w_7,7'b0};
assign c[1655:1472] = {84'b0,c_w_8,8'b0};
assign c[1839:1656] = {83'b0,c_w_9,9'b0};
assign c[2023:1840] = {82'b0,c_w_10,10'b0};
assign c[2207:2024] = {81'b0,c_w_11,11'b0};
assign c[2391:2208] = {80'b0,c_w_12,12'b0};
assign c[2575:2392] = {79'b0,c_w_13,13'b0};
assign c[2759:2576] = {78'b0,c_w_14,14'b0};
assign c[2943:2760] = {77'b0,c_w_15,15'b0};
assign c[3127:2944] = {76'b0,c_w_16,16'b0};
assign c[3311:3128] = {75'b0,c_w_17,17'b0};
assign c[3495:3312] = {74'b0,c_w_18,18'b0};
assign c[3679:3496] = {73'b0,c_w_19,19'b0};
assign c[3863:3680] = {72'b0,c_w_20,20'b0};
assign c[4047:3864] = {71'b0,c_w_21,21'b0};
assign c[4231:4048] = {70'b0,c_w_22,22'b0};
assign c[4415:4232] = {69'b0,c_w_23,23'b0};
assign c[4599:4416] = {68'b0,c_w_24,24'b0};
assign c[4783:4600] = {67'b0,c_w_25,25'b0};
assign c[4967:4784] = {66'b0,c_w_26,26'b0};
assign c[5151:4968] = {65'b0,c_w_27,27'b0};
assign c[5335:5152] = {64'b0,c_w_28,28'b0};
assign c[5519:5336] = {63'b0,c_w_29,29'b0};
assign c[5703:5520] = {62'b0,c_w_30,30'b0};
assign c[5887:5704] = {61'b0,c_w_31,31'b0};
assign c[6071:5888] = {60'b0,c_w_32,32'b0};
assign c[6255:6072] = {59'b0,c_w_33,33'b0};
assign c[6439:6256] = {58'b0,c_w_34,34'b0};
assign c[6623:6440] = {57'b0,c_w_35,35'b0};
assign c[6807:6624] = {56'b0,c_w_36,36'b0};
assign c[6991:6808] = {55'b0,c_w_37,37'b0};
assign c[7175:6992] = {54'b0,c_w_38,38'b0};
assign c[7359:7176] = {53'b0,c_w_39,39'b0};
assign c[7543:7360] = {52'b0,c_w_40,40'b0};
assign c[7727:7544] = {51'b0,c_w_41,41'b0};
assign c[7911:7728] = {50'b0,c_w_42,42'b0};
assign c[8095:7912] = {49'b0,c_w_43,43'b0};
assign c[8279:8096] = {48'b0,c_w_44,44'b0};
assign c[8463:8280] = {47'b0,c_w_45,45'b0};
assign c[8647:8464] = {46'b0,c_w_46,46'b0};
assign c[8831:8648] = {45'b0,c_w_47,47'b0};
assign c[9015:8832] = {44'b0,c_w_48,48'b0};
assign c[9199:9016] = {43'b0,c_w_49,49'b0};
assign c[9383:9200] = {42'b0,c_w_50,50'b0};
assign c[9567:9384] = {41'b0,c_w_51,51'b0};
assign c[9751:9568] = {40'b0,c_w_52,52'b0};
assign c[9935:9752] = {39'b0,c_w_53,53'b0};
assign c[10119:9936] = {38'b0,c_w_54,54'b0};
assign c[10303:10120] = {37'b0,c_w_55,55'b0};
assign c[10487:10304] = {36'b0,c_w_56,56'b0};
assign c[10671:10488] = {35'b0,c_w_57,57'b0};
assign c[10855:10672] = {34'b0,c_w_58,58'b0};
assign c[11039:10856] = {33'b0,c_w_59,59'b0};
assign c[11223:11040] = {32'b0,c_w_60,60'b0};
assign c[11407:11224] = {31'b0,c_w_61,61'b0};
assign c[11591:11408] = {30'b0,c_w_62,62'b0};
assign c[11775:11592] = {29'b0,c_w_63,63'b0};
assign c[11959:11776] = {28'b0,c_w_64,64'b0};
assign c[12143:11960] = {27'b0,c_w_65,65'b0};
assign c[12327:12144] = {26'b0,c_w_66,66'b0};
assign c[12511:12328] = {25'b0,c_w_67,67'b0};
assign c[12695:12512] = {24'b0,c_w_68,68'b0};
assign c[12879:12696] = {23'b0,c_w_69,69'b0};
assign c[13063:12880] = {22'b0,c_w_70,70'b0};
assign c[13247:13064] = {21'b0,c_w_71,71'b0};
assign c[13431:13248] = {20'b0,c_w_72,72'b0};
assign c[13615:13432] = {19'b0,c_w_73,73'b0};
assign c[13799:13616] = {18'b0,c_w_74,74'b0};
assign c[13983:13800] = {17'b0,c_w_75,75'b0};
assign c[14167:13984] = {16'b0,c_w_76,76'b0};
assign c[14351:14168] = {15'b0,c_w_77,77'b0};
assign c[14535:14352] = {14'b0,c_w_78,78'b0};
assign c[14719:14536] = {13'b0,c_w_79,79'b0};
assign c[14903:14720] = {12'b0,c_w_80,80'b0};
assign c[15087:14904] = {11'b0,c_w_81,81'b0};
assign c[15271:15088] = {10'b0,c_w_82,82'b0};
assign c[15455:15272] = {9'b0,c_w_83,83'b0};
assign c[15639:15456] = {8'b0,c_w_84,84'b0};
assign c[15823:15640] = {7'b0,c_w_85,85'b0};
assign c[16007:15824] = {6'b0,c_w_86,86'b0};
assign c[16191:16008] = {5'b0,c_w_87,87'b0};
assign c[16375:16192] = {4'b0,c_w_88,88'b0};
assign c[16559:16376] = {3'b0,c_w_89,89'b0};
assign c[16743:16560] = {2'b0,c_w_90,90'b0};
assign c[16927:16744] = {1'b0,c_w_91,91'b0};
    
endmodule
    