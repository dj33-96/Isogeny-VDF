

module csa_tree_92x184(
    input [16927:0] A, // lines are appended together
    output[183:0] B_0,
    output[183:0] B_1
);

wire [11407:0] tree_1;
wire [7727:0] tree_2;
wire [5151:0] tree_3;
wire [3495:0] tree_4;
wire [2391:0] tree_5;
wire [1655:0] tree_6;
wire [1103:0] tree_7;
wire [735:0] tree_8;
wire [551:0] tree_9;
wire [367:0] tree_10;
// layer-1
csa_184 csau_184_i0(A[183:0],A[367:184],A[551:368],tree_1[183:0],tree_1[367:184]);
csa_184 csau_184_i1(A[735:552],A[919:736],A[1103:920],tree_1[551:368],tree_1[735:552]);
csa_184 csau_184_i2(A[1287:1104],A[1471:1288],A[1655:1472],tree_1[919:736],tree_1[1103:920]);
csa_184 csau_184_i3(A[1839:1656],A[2023:1840],A[2207:2024],tree_1[1287:1104],tree_1[1471:1288]);
csa_184 csau_184_i4(A[2391:2208],A[2575:2392],A[2759:2576],tree_1[1655:1472],tree_1[1839:1656]);
csa_184 csau_184_i5(A[2943:2760],A[3127:2944],A[3311:3128],tree_1[2023:1840],tree_1[2207:2024]);
csa_184 csau_184_i6(A[3495:3312],A[3679:3496],A[3863:3680],tree_1[2391:2208],tree_1[2575:2392]);
csa_184 csau_184_i7(A[4047:3864],A[4231:4048],A[4415:4232],tree_1[2759:2576],tree_1[2943:2760]);
csa_184 csau_184_i8(A[4599:4416],A[4783:4600],A[4967:4784],tree_1[3127:2944],tree_1[3311:3128]);
csa_184 csau_184_i9(A[5151:4968],A[5335:5152],A[5519:5336],tree_1[3495:3312],tree_1[3679:3496]);
csa_184 csau_184_i10(A[5703:5520],A[5887:5704],A[6071:5888],tree_1[3863:3680],tree_1[4047:3864]);
csa_184 csau_184_i11(A[6255:6072],A[6439:6256],A[6623:6440],tree_1[4231:4048],tree_1[4415:4232]);
csa_184 csau_184_i12(A[6807:6624],A[6991:6808],A[7175:6992],tree_1[4599:4416],tree_1[4783:4600]);
csa_184 csau_184_i13(A[7359:7176],A[7543:7360],A[7727:7544],tree_1[4967:4784],tree_1[5151:4968]);
csa_184 csau_184_i14(A[7911:7728],A[8095:7912],A[8279:8096],tree_1[5335:5152],tree_1[5519:5336]);
csa_184 csau_184_i15(A[8463:8280],A[8647:8464],A[8831:8648],tree_1[5703:5520],tree_1[5887:5704]);
csa_184 csau_184_i16(A[9015:8832],A[9199:9016],A[9383:9200],tree_1[6071:5888],tree_1[6255:6072]);
csa_184 csau_184_i17(A[9567:9384],A[9751:9568],A[9935:9752],tree_1[6439:6256],tree_1[6623:6440]);
csa_184 csau_184_i18(A[10119:9936],A[10303:10120],A[10487:10304],tree_1[6807:6624],tree_1[6991:6808]);
csa_184 csau_184_i19(A[10671:10488],A[10855:10672],A[11039:10856],tree_1[7175:6992],tree_1[7359:7176]);
csa_184 csau_184_i20(A[11223:11040],A[11407:11224],A[11591:11408],tree_1[7543:7360],tree_1[7727:7544]);
csa_184 csau_184_i21(A[11775:11592],A[11959:11776],A[12143:11960],tree_1[7911:7728],tree_1[8095:7912]);
csa_184 csau_184_i22(A[12327:12144],A[12511:12328],A[12695:12512],tree_1[8279:8096],tree_1[8463:8280]);
csa_184 csau_184_i23(A[12879:12696],A[13063:12880],A[13247:13064],tree_1[8647:8464],tree_1[8831:8648]);
csa_184 csau_184_i24(A[13431:13248],A[13615:13432],A[13799:13616],tree_1[9015:8832],tree_1[9199:9016]);
csa_184 csau_184_i25(A[13983:13800],A[14167:13984],A[14351:14168],tree_1[9383:9200],tree_1[9567:9384]);
csa_184 csau_184_i26(A[14535:14352],A[14719:14536],A[14903:14720],tree_1[9751:9568],tree_1[9935:9752]);
csa_184 csau_184_i27(A[15087:14904],A[15271:15088],A[15455:15272],tree_1[10119:9936],tree_1[10303:10120]);
csa_184 csau_184_i28(A[15639:15456],A[15823:15640],A[16007:15824],tree_1[10487:10304],tree_1[10671:10488]);
csa_184 csau_184_i29(A[16191:16008],A[16375:16192],A[16559:16376],tree_1[10855:10672],tree_1[11039:10856]);
assign tree_1[11223:11040] = A[16743:16560];
assign tree_1[11407:11224] = A[16927:16744];
// layer-2
csa_184 csau_184_i30(tree_1[183:0],tree_1[367:184],tree_1[551:368],tree_2[183:0],tree_2[367:184]);
csa_184 csau_184_i31(tree_1[735:552],tree_1[919:736],tree_1[1103:920],tree_2[551:368],tree_2[735:552]);
csa_184 csau_184_i32(tree_1[1287:1104],tree_1[1471:1288],tree_1[1655:1472],tree_2[919:736],tree_2[1103:920]);
csa_184 csau_184_i33(tree_1[1839:1656],tree_1[2023:1840],tree_1[2207:2024],tree_2[1287:1104],tree_2[1471:1288]);
csa_184 csau_184_i34(tree_1[2391:2208],tree_1[2575:2392],tree_1[2759:2576],tree_2[1655:1472],tree_2[1839:1656]);
csa_184 csau_184_i35(tree_1[2943:2760],tree_1[3127:2944],tree_1[3311:3128],tree_2[2023:1840],tree_2[2207:2024]);
csa_184 csau_184_i36(tree_1[3495:3312],tree_1[3679:3496],tree_1[3863:3680],tree_2[2391:2208],tree_2[2575:2392]);
csa_184 csau_184_i37(tree_1[4047:3864],tree_1[4231:4048],tree_1[4415:4232],tree_2[2759:2576],tree_2[2943:2760]);
csa_184 csau_184_i38(tree_1[4599:4416],tree_1[4783:4600],tree_1[4967:4784],tree_2[3127:2944],tree_2[3311:3128]);
csa_184 csau_184_i39(tree_1[5151:4968],tree_1[5335:5152],tree_1[5519:5336],tree_2[3495:3312],tree_2[3679:3496]);
csa_184 csau_184_i40(tree_1[5703:5520],tree_1[5887:5704],tree_1[6071:5888],tree_2[3863:3680],tree_2[4047:3864]);
csa_184 csau_184_i41(tree_1[6255:6072],tree_1[6439:6256],tree_1[6623:6440],tree_2[4231:4048],tree_2[4415:4232]);
csa_184 csau_184_i42(tree_1[6807:6624],tree_1[6991:6808],tree_1[7175:6992],tree_2[4599:4416],tree_2[4783:4600]);
csa_184 csau_184_i43(tree_1[7359:7176],tree_1[7543:7360],tree_1[7727:7544],tree_2[4967:4784],tree_2[5151:4968]);
csa_184 csau_184_i44(tree_1[7911:7728],tree_1[8095:7912],tree_1[8279:8096],tree_2[5335:5152],tree_2[5519:5336]);
csa_184 csau_184_i45(tree_1[8463:8280],tree_1[8647:8464],tree_1[8831:8648],tree_2[5703:5520],tree_2[5887:5704]);
csa_184 csau_184_i46(tree_1[9015:8832],tree_1[9199:9016],tree_1[9383:9200],tree_2[6071:5888],tree_2[6255:6072]);
csa_184 csau_184_i47(tree_1[9567:9384],tree_1[9751:9568],tree_1[9935:9752],tree_2[6439:6256],tree_2[6623:6440]);
csa_184 csau_184_i48(tree_1[10119:9936],tree_1[10303:10120],tree_1[10487:10304],tree_2[6807:6624],tree_2[6991:6808]);
csa_184 csau_184_i49(tree_1[10671:10488],tree_1[10855:10672],tree_1[11039:10856],tree_2[7175:6992],tree_2[7359:7176]);
assign tree_2[7543:7360] = tree_1[11223:11040];
assign tree_2[7727:7544] = tree_1[11407:11224];
// layer-3
csa_184 csau_184_i50(tree_2[183:0],tree_2[367:184],tree_2[551:368],tree_3[183:0],tree_3[367:184]);
csa_184 csau_184_i51(tree_2[735:552],tree_2[919:736],tree_2[1103:920],tree_3[551:368],tree_3[735:552]);
csa_184 csau_184_i52(tree_2[1287:1104],tree_2[1471:1288],tree_2[1655:1472],tree_3[919:736],tree_3[1103:920]);
csa_184 csau_184_i53(tree_2[1839:1656],tree_2[2023:1840],tree_2[2207:2024],tree_3[1287:1104],tree_3[1471:1288]);
csa_184 csau_184_i54(tree_2[2391:2208],tree_2[2575:2392],tree_2[2759:2576],tree_3[1655:1472],tree_3[1839:1656]);
csa_184 csau_184_i55(tree_2[2943:2760],tree_2[3127:2944],tree_2[3311:3128],tree_3[2023:1840],tree_3[2207:2024]);
csa_184 csau_184_i56(tree_2[3495:3312],tree_2[3679:3496],tree_2[3863:3680],tree_3[2391:2208],tree_3[2575:2392]);
csa_184 csau_184_i57(tree_2[4047:3864],tree_2[4231:4048],tree_2[4415:4232],tree_3[2759:2576],tree_3[2943:2760]);
csa_184 csau_184_i58(tree_2[4599:4416],tree_2[4783:4600],tree_2[4967:4784],tree_3[3127:2944],tree_3[3311:3128]);
csa_184 csau_184_i59(tree_2[5151:4968],tree_2[5335:5152],tree_2[5519:5336],tree_3[3495:3312],tree_3[3679:3496]);
csa_184 csau_184_i60(tree_2[5703:5520],tree_2[5887:5704],tree_2[6071:5888],tree_3[3863:3680],tree_3[4047:3864]);
csa_184 csau_184_i61(tree_2[6255:6072],tree_2[6439:6256],tree_2[6623:6440],tree_3[4231:4048],tree_3[4415:4232]);
csa_184 csau_184_i62(tree_2[6807:6624],tree_2[6991:6808],tree_2[7175:6992],tree_3[4599:4416],tree_3[4783:4600]);
csa_184 csau_184_i63(tree_2[7359:7176],tree_2[7543:7360],tree_2[7727:7544],tree_3[4967:4784],tree_3[5151:4968]);
// layer-4
csa_184 csau_184_i64(tree_3[183:0],tree_3[367:184],tree_3[551:368],tree_4[183:0],tree_4[367:184]);
csa_184 csau_184_i65(tree_3[735:552],tree_3[919:736],tree_3[1103:920],tree_4[551:368],tree_4[735:552]);
csa_184 csau_184_i66(tree_3[1287:1104],tree_3[1471:1288],tree_3[1655:1472],tree_4[919:736],tree_4[1103:920]);
csa_184 csau_184_i67(tree_3[1839:1656],tree_3[2023:1840],tree_3[2207:2024],tree_4[1287:1104],tree_4[1471:1288]);
csa_184 csau_184_i68(tree_3[2391:2208],tree_3[2575:2392],tree_3[2759:2576],tree_4[1655:1472],tree_4[1839:1656]);
csa_184 csau_184_i69(tree_3[2943:2760],tree_3[3127:2944],tree_3[3311:3128],tree_4[2023:1840],tree_4[2207:2024]);
csa_184 csau_184_i70(tree_3[3495:3312],tree_3[3679:3496],tree_3[3863:3680],tree_4[2391:2208],tree_4[2575:2392]);
csa_184 csau_184_i71(tree_3[4047:3864],tree_3[4231:4048],tree_3[4415:4232],tree_4[2759:2576],tree_4[2943:2760]);
csa_184 csau_184_i72(tree_3[4599:4416],tree_3[4783:4600],tree_3[4967:4784],tree_4[3127:2944],tree_4[3311:3128]);
assign tree_4[3495:3312] = tree_3[5151:4968];
// layer-5
csa_184 csau_184_i73(tree_4[183:0],tree_4[367:184],tree_4[551:368],tree_5[183:0],tree_5[367:184]);
csa_184 csau_184_i74(tree_4[735:552],tree_4[919:736],tree_4[1103:920],tree_5[551:368],tree_5[735:552]);
csa_184 csau_184_i75(tree_4[1287:1104],tree_4[1471:1288],tree_4[1655:1472],tree_5[919:736],tree_5[1103:920]);
csa_184 csau_184_i76(tree_4[1839:1656],tree_4[2023:1840],tree_4[2207:2024],tree_5[1287:1104],tree_5[1471:1288]);
csa_184 csau_184_i77(tree_4[2391:2208],tree_4[2575:2392],tree_4[2759:2576],tree_5[1655:1472],tree_5[1839:1656]);
csa_184 csau_184_i78(tree_4[2943:2760],tree_4[3127:2944],tree_4[3311:3128],tree_5[2023:1840],tree_5[2207:2024]);
assign tree_5[2391:2208] = tree_4[3495:3312];
// layer-6
csa_184 csau_184_i79(tree_5[183:0],tree_5[367:184],tree_5[551:368],tree_6[183:0],tree_6[367:184]);
csa_184 csau_184_i80(tree_5[735:552],tree_5[919:736],tree_5[1103:920],tree_6[551:368],tree_6[735:552]);
csa_184 csau_184_i81(tree_5[1287:1104],tree_5[1471:1288],tree_5[1655:1472],tree_6[919:736],tree_6[1103:920]);
csa_184 csau_184_i82(tree_5[1839:1656],tree_5[2023:1840],tree_5[2207:2024],tree_6[1287:1104],tree_6[1471:1288]);
assign tree_6[1655:1472] = tree_5[2391:2208];
// layer-7
csa_184 csau_184_i83(tree_6[183:0],tree_6[367:184],tree_6[551:368],tree_7[183:0],tree_7[367:184]);
csa_184 csau_184_i84(tree_6[735:552],tree_6[919:736],tree_6[1103:920],tree_7[551:368],tree_7[735:552]);
csa_184 csau_184_i85(tree_6[1287:1104],tree_6[1471:1288],tree_6[1655:1472],tree_7[919:736],tree_7[1103:920]);
// layer-8
csa_184 csau_184_i86(tree_7[183:0],tree_7[367:184],tree_7[551:368],tree_8[183:0],tree_8[367:184]);
csa_184 csau_184_i87(tree_7[735:552],tree_7[919:736],tree_7[1103:920],tree_8[551:368],tree_8[735:552]);
// layer-9
csa_184 csau_184_i88(tree_8[183:0],tree_8[367:184],tree_8[551:368],tree_9[183:0],tree_9[367:184]);
assign tree_9[551:368] = tree_8[735:552];
// layer-10
csa_184 csau_184_i89(tree_9[183:0],tree_9[367:184],tree_9[551:368],tree_10[183:0],tree_10[367:184]);

// final assignment
assign B_0 = tree_10[183:0];
assign B_1 = tree_10[367:184];

endmodule
