
module xor_89_array(
    input [88:0] in0,in1,
    output [88:0] out0
);

assign out0 = in0 ^ in1;

endmodule
    