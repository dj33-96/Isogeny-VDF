

module csa_tree_1509x3018(
    input [4554161:0] A, // lines are appended together
    output[3017:0] B_0,
    output[3017:0] B_1
);

wire [3036107:0] tree_1;
wire [2025077:0] tree_2;
wire [1352063:0] tree_3;
wire [902381:0] tree_4;
wire [603599:0] tree_5;
wire [404411:0] tree_6;
wire [271619:0] tree_7;
wire [181079:0] tree_8;
wire [120719:0] tree_9;
wire [81485:0] tree_10;
wire [54323:0] tree_11;
wire [36215:0] tree_12;
wire [24143:0] tree_13;
wire [18107:0] tree_14;
wire [12071:0] tree_15;
wire [9053:0] tree_16;
wire [6035:0] tree_17;
// layer-1
csa_3018 csau_3018_i0(A[3017:0],A[6035:3018],A[9053:6036],tree_1[3017:0],tree_1[6035:3018]);
csa_3018 csau_3018_i1(A[12071:9054],A[15089:12072],A[18107:15090],tree_1[9053:6036],tree_1[12071:9054]);
csa_3018 csau_3018_i2(A[21125:18108],A[24143:21126],A[27161:24144],tree_1[15089:12072],tree_1[18107:15090]);
csa_3018 csau_3018_i3(A[30179:27162],A[33197:30180],A[36215:33198],tree_1[21125:18108],tree_1[24143:21126]);
csa_3018 csau_3018_i4(A[39233:36216],A[42251:39234],A[45269:42252],tree_1[27161:24144],tree_1[30179:27162]);
csa_3018 csau_3018_i5(A[48287:45270],A[51305:48288],A[54323:51306],tree_1[33197:30180],tree_1[36215:33198]);
csa_3018 csau_3018_i6(A[57341:54324],A[60359:57342],A[63377:60360],tree_1[39233:36216],tree_1[42251:39234]);
csa_3018 csau_3018_i7(A[66395:63378],A[69413:66396],A[72431:69414],tree_1[45269:42252],tree_1[48287:45270]);
csa_3018 csau_3018_i8(A[75449:72432],A[78467:75450],A[81485:78468],tree_1[51305:48288],tree_1[54323:51306]);
csa_3018 csau_3018_i9(A[84503:81486],A[87521:84504],A[90539:87522],tree_1[57341:54324],tree_1[60359:57342]);
csa_3018 csau_3018_i10(A[93557:90540],A[96575:93558],A[99593:96576],tree_1[63377:60360],tree_1[66395:63378]);
csa_3018 csau_3018_i11(A[102611:99594],A[105629:102612],A[108647:105630],tree_1[69413:66396],tree_1[72431:69414]);
csa_3018 csau_3018_i12(A[111665:108648],A[114683:111666],A[117701:114684],tree_1[75449:72432],tree_1[78467:75450]);
csa_3018 csau_3018_i13(A[120719:117702],A[123737:120720],A[126755:123738],tree_1[81485:78468],tree_1[84503:81486]);
csa_3018 csau_3018_i14(A[129773:126756],A[132791:129774],A[135809:132792],tree_1[87521:84504],tree_1[90539:87522]);
csa_3018 csau_3018_i15(A[138827:135810],A[141845:138828],A[144863:141846],tree_1[93557:90540],tree_1[96575:93558]);
csa_3018 csau_3018_i16(A[147881:144864],A[150899:147882],A[153917:150900],tree_1[99593:96576],tree_1[102611:99594]);
csa_3018 csau_3018_i17(A[156935:153918],A[159953:156936],A[162971:159954],tree_1[105629:102612],tree_1[108647:105630]);
csa_3018 csau_3018_i18(A[165989:162972],A[169007:165990],A[172025:169008],tree_1[111665:108648],tree_1[114683:111666]);
csa_3018 csau_3018_i19(A[175043:172026],A[178061:175044],A[181079:178062],tree_1[117701:114684],tree_1[120719:117702]);
csa_3018 csau_3018_i20(A[184097:181080],A[187115:184098],A[190133:187116],tree_1[123737:120720],tree_1[126755:123738]);
csa_3018 csau_3018_i21(A[193151:190134],A[196169:193152],A[199187:196170],tree_1[129773:126756],tree_1[132791:129774]);
csa_3018 csau_3018_i22(A[202205:199188],A[205223:202206],A[208241:205224],tree_1[135809:132792],tree_1[138827:135810]);
csa_3018 csau_3018_i23(A[211259:208242],A[214277:211260],A[217295:214278],tree_1[141845:138828],tree_1[144863:141846]);
csa_3018 csau_3018_i24(A[220313:217296],A[223331:220314],A[226349:223332],tree_1[147881:144864],tree_1[150899:147882]);
csa_3018 csau_3018_i25(A[229367:226350],A[232385:229368],A[235403:232386],tree_1[153917:150900],tree_1[156935:153918]);
csa_3018 csau_3018_i26(A[238421:235404],A[241439:238422],A[244457:241440],tree_1[159953:156936],tree_1[162971:159954]);
csa_3018 csau_3018_i27(A[247475:244458],A[250493:247476],A[253511:250494],tree_1[165989:162972],tree_1[169007:165990]);
csa_3018 csau_3018_i28(A[256529:253512],A[259547:256530],A[262565:259548],tree_1[172025:169008],tree_1[175043:172026]);
csa_3018 csau_3018_i29(A[265583:262566],A[268601:265584],A[271619:268602],tree_1[178061:175044],tree_1[181079:178062]);
csa_3018 csau_3018_i30(A[274637:271620],A[277655:274638],A[280673:277656],tree_1[184097:181080],tree_1[187115:184098]);
csa_3018 csau_3018_i31(A[283691:280674],A[286709:283692],A[289727:286710],tree_1[190133:187116],tree_1[193151:190134]);
csa_3018 csau_3018_i32(A[292745:289728],A[295763:292746],A[298781:295764],tree_1[196169:193152],tree_1[199187:196170]);
csa_3018 csau_3018_i33(A[301799:298782],A[304817:301800],A[307835:304818],tree_1[202205:199188],tree_1[205223:202206]);
csa_3018 csau_3018_i34(A[310853:307836],A[313871:310854],A[316889:313872],tree_1[208241:205224],tree_1[211259:208242]);
csa_3018 csau_3018_i35(A[319907:316890],A[322925:319908],A[325943:322926],tree_1[214277:211260],tree_1[217295:214278]);
csa_3018 csau_3018_i36(A[328961:325944],A[331979:328962],A[334997:331980],tree_1[220313:217296],tree_1[223331:220314]);
csa_3018 csau_3018_i37(A[338015:334998],A[341033:338016],A[344051:341034],tree_1[226349:223332],tree_1[229367:226350]);
csa_3018 csau_3018_i38(A[347069:344052],A[350087:347070],A[353105:350088],tree_1[232385:229368],tree_1[235403:232386]);
csa_3018 csau_3018_i39(A[356123:353106],A[359141:356124],A[362159:359142],tree_1[238421:235404],tree_1[241439:238422]);
csa_3018 csau_3018_i40(A[365177:362160],A[368195:365178],A[371213:368196],tree_1[244457:241440],tree_1[247475:244458]);
csa_3018 csau_3018_i41(A[374231:371214],A[377249:374232],A[380267:377250],tree_1[250493:247476],tree_1[253511:250494]);
csa_3018 csau_3018_i42(A[383285:380268],A[386303:383286],A[389321:386304],tree_1[256529:253512],tree_1[259547:256530]);
csa_3018 csau_3018_i43(A[392339:389322],A[395357:392340],A[398375:395358],tree_1[262565:259548],tree_1[265583:262566]);
csa_3018 csau_3018_i44(A[401393:398376],A[404411:401394],A[407429:404412],tree_1[268601:265584],tree_1[271619:268602]);
csa_3018 csau_3018_i45(A[410447:407430],A[413465:410448],A[416483:413466],tree_1[274637:271620],tree_1[277655:274638]);
csa_3018 csau_3018_i46(A[419501:416484],A[422519:419502],A[425537:422520],tree_1[280673:277656],tree_1[283691:280674]);
csa_3018 csau_3018_i47(A[428555:425538],A[431573:428556],A[434591:431574],tree_1[286709:283692],tree_1[289727:286710]);
csa_3018 csau_3018_i48(A[437609:434592],A[440627:437610],A[443645:440628],tree_1[292745:289728],tree_1[295763:292746]);
csa_3018 csau_3018_i49(A[446663:443646],A[449681:446664],A[452699:449682],tree_1[298781:295764],tree_1[301799:298782]);
csa_3018 csau_3018_i50(A[455717:452700],A[458735:455718],A[461753:458736],tree_1[304817:301800],tree_1[307835:304818]);
csa_3018 csau_3018_i51(A[464771:461754],A[467789:464772],A[470807:467790],tree_1[310853:307836],tree_1[313871:310854]);
csa_3018 csau_3018_i52(A[473825:470808],A[476843:473826],A[479861:476844],tree_1[316889:313872],tree_1[319907:316890]);
csa_3018 csau_3018_i53(A[482879:479862],A[485897:482880],A[488915:485898],tree_1[322925:319908],tree_1[325943:322926]);
csa_3018 csau_3018_i54(A[491933:488916],A[494951:491934],A[497969:494952],tree_1[328961:325944],tree_1[331979:328962]);
csa_3018 csau_3018_i55(A[500987:497970],A[504005:500988],A[507023:504006],tree_1[334997:331980],tree_1[338015:334998]);
csa_3018 csau_3018_i56(A[510041:507024],A[513059:510042],A[516077:513060],tree_1[341033:338016],tree_1[344051:341034]);
csa_3018 csau_3018_i57(A[519095:516078],A[522113:519096],A[525131:522114],tree_1[347069:344052],tree_1[350087:347070]);
csa_3018 csau_3018_i58(A[528149:525132],A[531167:528150],A[534185:531168],tree_1[353105:350088],tree_1[356123:353106]);
csa_3018 csau_3018_i59(A[537203:534186],A[540221:537204],A[543239:540222],tree_1[359141:356124],tree_1[362159:359142]);
csa_3018 csau_3018_i60(A[546257:543240],A[549275:546258],A[552293:549276],tree_1[365177:362160],tree_1[368195:365178]);
csa_3018 csau_3018_i61(A[555311:552294],A[558329:555312],A[561347:558330],tree_1[371213:368196],tree_1[374231:371214]);
csa_3018 csau_3018_i62(A[564365:561348],A[567383:564366],A[570401:567384],tree_1[377249:374232],tree_1[380267:377250]);
csa_3018 csau_3018_i63(A[573419:570402],A[576437:573420],A[579455:576438],tree_1[383285:380268],tree_1[386303:383286]);
csa_3018 csau_3018_i64(A[582473:579456],A[585491:582474],A[588509:585492],tree_1[389321:386304],tree_1[392339:389322]);
csa_3018 csau_3018_i65(A[591527:588510],A[594545:591528],A[597563:594546],tree_1[395357:392340],tree_1[398375:395358]);
csa_3018 csau_3018_i66(A[600581:597564],A[603599:600582],A[606617:603600],tree_1[401393:398376],tree_1[404411:401394]);
csa_3018 csau_3018_i67(A[609635:606618],A[612653:609636],A[615671:612654],tree_1[407429:404412],tree_1[410447:407430]);
csa_3018 csau_3018_i68(A[618689:615672],A[621707:618690],A[624725:621708],tree_1[413465:410448],tree_1[416483:413466]);
csa_3018 csau_3018_i69(A[627743:624726],A[630761:627744],A[633779:630762],tree_1[419501:416484],tree_1[422519:419502]);
csa_3018 csau_3018_i70(A[636797:633780],A[639815:636798],A[642833:639816],tree_1[425537:422520],tree_1[428555:425538]);
csa_3018 csau_3018_i71(A[645851:642834],A[648869:645852],A[651887:648870],tree_1[431573:428556],tree_1[434591:431574]);
csa_3018 csau_3018_i72(A[654905:651888],A[657923:654906],A[660941:657924],tree_1[437609:434592],tree_1[440627:437610]);
csa_3018 csau_3018_i73(A[663959:660942],A[666977:663960],A[669995:666978],tree_1[443645:440628],tree_1[446663:443646]);
csa_3018 csau_3018_i74(A[673013:669996],A[676031:673014],A[679049:676032],tree_1[449681:446664],tree_1[452699:449682]);
csa_3018 csau_3018_i75(A[682067:679050],A[685085:682068],A[688103:685086],tree_1[455717:452700],tree_1[458735:455718]);
csa_3018 csau_3018_i76(A[691121:688104],A[694139:691122],A[697157:694140],tree_1[461753:458736],tree_1[464771:461754]);
csa_3018 csau_3018_i77(A[700175:697158],A[703193:700176],A[706211:703194],tree_1[467789:464772],tree_1[470807:467790]);
csa_3018 csau_3018_i78(A[709229:706212],A[712247:709230],A[715265:712248],tree_1[473825:470808],tree_1[476843:473826]);
csa_3018 csau_3018_i79(A[718283:715266],A[721301:718284],A[724319:721302],tree_1[479861:476844],tree_1[482879:479862]);
csa_3018 csau_3018_i80(A[727337:724320],A[730355:727338],A[733373:730356],tree_1[485897:482880],tree_1[488915:485898]);
csa_3018 csau_3018_i81(A[736391:733374],A[739409:736392],A[742427:739410],tree_1[491933:488916],tree_1[494951:491934]);
csa_3018 csau_3018_i82(A[745445:742428],A[748463:745446],A[751481:748464],tree_1[497969:494952],tree_1[500987:497970]);
csa_3018 csau_3018_i83(A[754499:751482],A[757517:754500],A[760535:757518],tree_1[504005:500988],tree_1[507023:504006]);
csa_3018 csau_3018_i84(A[763553:760536],A[766571:763554],A[769589:766572],tree_1[510041:507024],tree_1[513059:510042]);
csa_3018 csau_3018_i85(A[772607:769590],A[775625:772608],A[778643:775626],tree_1[516077:513060],tree_1[519095:516078]);
csa_3018 csau_3018_i86(A[781661:778644],A[784679:781662],A[787697:784680],tree_1[522113:519096],tree_1[525131:522114]);
csa_3018 csau_3018_i87(A[790715:787698],A[793733:790716],A[796751:793734],tree_1[528149:525132],tree_1[531167:528150]);
csa_3018 csau_3018_i88(A[799769:796752],A[802787:799770],A[805805:802788],tree_1[534185:531168],tree_1[537203:534186]);
csa_3018 csau_3018_i89(A[808823:805806],A[811841:808824],A[814859:811842],tree_1[540221:537204],tree_1[543239:540222]);
csa_3018 csau_3018_i90(A[817877:814860],A[820895:817878],A[823913:820896],tree_1[546257:543240],tree_1[549275:546258]);
csa_3018 csau_3018_i91(A[826931:823914],A[829949:826932],A[832967:829950],tree_1[552293:549276],tree_1[555311:552294]);
csa_3018 csau_3018_i92(A[835985:832968],A[839003:835986],A[842021:839004],tree_1[558329:555312],tree_1[561347:558330]);
csa_3018 csau_3018_i93(A[845039:842022],A[848057:845040],A[851075:848058],tree_1[564365:561348],tree_1[567383:564366]);
csa_3018 csau_3018_i94(A[854093:851076],A[857111:854094],A[860129:857112],tree_1[570401:567384],tree_1[573419:570402]);
csa_3018 csau_3018_i95(A[863147:860130],A[866165:863148],A[869183:866166],tree_1[576437:573420],tree_1[579455:576438]);
csa_3018 csau_3018_i96(A[872201:869184],A[875219:872202],A[878237:875220],tree_1[582473:579456],tree_1[585491:582474]);
csa_3018 csau_3018_i97(A[881255:878238],A[884273:881256],A[887291:884274],tree_1[588509:585492],tree_1[591527:588510]);
csa_3018 csau_3018_i98(A[890309:887292],A[893327:890310],A[896345:893328],tree_1[594545:591528],tree_1[597563:594546]);
csa_3018 csau_3018_i99(A[899363:896346],A[902381:899364],A[905399:902382],tree_1[600581:597564],tree_1[603599:600582]);
csa_3018 csau_3018_i100(A[908417:905400],A[911435:908418],A[914453:911436],tree_1[606617:603600],tree_1[609635:606618]);
csa_3018 csau_3018_i101(A[917471:914454],A[920489:917472],A[923507:920490],tree_1[612653:609636],tree_1[615671:612654]);
csa_3018 csau_3018_i102(A[926525:923508],A[929543:926526],A[932561:929544],tree_1[618689:615672],tree_1[621707:618690]);
csa_3018 csau_3018_i103(A[935579:932562],A[938597:935580],A[941615:938598],tree_1[624725:621708],tree_1[627743:624726]);
csa_3018 csau_3018_i104(A[944633:941616],A[947651:944634],A[950669:947652],tree_1[630761:627744],tree_1[633779:630762]);
csa_3018 csau_3018_i105(A[953687:950670],A[956705:953688],A[959723:956706],tree_1[636797:633780],tree_1[639815:636798]);
csa_3018 csau_3018_i106(A[962741:959724],A[965759:962742],A[968777:965760],tree_1[642833:639816],tree_1[645851:642834]);
csa_3018 csau_3018_i107(A[971795:968778],A[974813:971796],A[977831:974814],tree_1[648869:645852],tree_1[651887:648870]);
csa_3018 csau_3018_i108(A[980849:977832],A[983867:980850],A[986885:983868],tree_1[654905:651888],tree_1[657923:654906]);
csa_3018 csau_3018_i109(A[989903:986886],A[992921:989904],A[995939:992922],tree_1[660941:657924],tree_1[663959:660942]);
csa_3018 csau_3018_i110(A[998957:995940],A[1001975:998958],A[1004993:1001976],tree_1[666977:663960],tree_1[669995:666978]);
csa_3018 csau_3018_i111(A[1008011:1004994],A[1011029:1008012],A[1014047:1011030],tree_1[673013:669996],tree_1[676031:673014]);
csa_3018 csau_3018_i112(A[1017065:1014048],A[1020083:1017066],A[1023101:1020084],tree_1[679049:676032],tree_1[682067:679050]);
csa_3018 csau_3018_i113(A[1026119:1023102],A[1029137:1026120],A[1032155:1029138],tree_1[685085:682068],tree_1[688103:685086]);
csa_3018 csau_3018_i114(A[1035173:1032156],A[1038191:1035174],A[1041209:1038192],tree_1[691121:688104],tree_1[694139:691122]);
csa_3018 csau_3018_i115(A[1044227:1041210],A[1047245:1044228],A[1050263:1047246],tree_1[697157:694140],tree_1[700175:697158]);
csa_3018 csau_3018_i116(A[1053281:1050264],A[1056299:1053282],A[1059317:1056300],tree_1[703193:700176],tree_1[706211:703194]);
csa_3018 csau_3018_i117(A[1062335:1059318],A[1065353:1062336],A[1068371:1065354],tree_1[709229:706212],tree_1[712247:709230]);
csa_3018 csau_3018_i118(A[1071389:1068372],A[1074407:1071390],A[1077425:1074408],tree_1[715265:712248],tree_1[718283:715266]);
csa_3018 csau_3018_i119(A[1080443:1077426],A[1083461:1080444],A[1086479:1083462],tree_1[721301:718284],tree_1[724319:721302]);
csa_3018 csau_3018_i120(A[1089497:1086480],A[1092515:1089498],A[1095533:1092516],tree_1[727337:724320],tree_1[730355:727338]);
csa_3018 csau_3018_i121(A[1098551:1095534],A[1101569:1098552],A[1104587:1101570],tree_1[733373:730356],tree_1[736391:733374]);
csa_3018 csau_3018_i122(A[1107605:1104588],A[1110623:1107606],A[1113641:1110624],tree_1[739409:736392],tree_1[742427:739410]);
csa_3018 csau_3018_i123(A[1116659:1113642],A[1119677:1116660],A[1122695:1119678],tree_1[745445:742428],tree_1[748463:745446]);
csa_3018 csau_3018_i124(A[1125713:1122696],A[1128731:1125714],A[1131749:1128732],tree_1[751481:748464],tree_1[754499:751482]);
csa_3018 csau_3018_i125(A[1134767:1131750],A[1137785:1134768],A[1140803:1137786],tree_1[757517:754500],tree_1[760535:757518]);
csa_3018 csau_3018_i126(A[1143821:1140804],A[1146839:1143822],A[1149857:1146840],tree_1[763553:760536],tree_1[766571:763554]);
csa_3018 csau_3018_i127(A[1152875:1149858],A[1155893:1152876],A[1158911:1155894],tree_1[769589:766572],tree_1[772607:769590]);
csa_3018 csau_3018_i128(A[1161929:1158912],A[1164947:1161930],A[1167965:1164948],tree_1[775625:772608],tree_1[778643:775626]);
csa_3018 csau_3018_i129(A[1170983:1167966],A[1174001:1170984],A[1177019:1174002],tree_1[781661:778644],tree_1[784679:781662]);
csa_3018 csau_3018_i130(A[1180037:1177020],A[1183055:1180038],A[1186073:1183056],tree_1[787697:784680],tree_1[790715:787698]);
csa_3018 csau_3018_i131(A[1189091:1186074],A[1192109:1189092],A[1195127:1192110],tree_1[793733:790716],tree_1[796751:793734]);
csa_3018 csau_3018_i132(A[1198145:1195128],A[1201163:1198146],A[1204181:1201164],tree_1[799769:796752],tree_1[802787:799770]);
csa_3018 csau_3018_i133(A[1207199:1204182],A[1210217:1207200],A[1213235:1210218],tree_1[805805:802788],tree_1[808823:805806]);
csa_3018 csau_3018_i134(A[1216253:1213236],A[1219271:1216254],A[1222289:1219272],tree_1[811841:808824],tree_1[814859:811842]);
csa_3018 csau_3018_i135(A[1225307:1222290],A[1228325:1225308],A[1231343:1228326],tree_1[817877:814860],tree_1[820895:817878]);
csa_3018 csau_3018_i136(A[1234361:1231344],A[1237379:1234362],A[1240397:1237380],tree_1[823913:820896],tree_1[826931:823914]);
csa_3018 csau_3018_i137(A[1243415:1240398],A[1246433:1243416],A[1249451:1246434],tree_1[829949:826932],tree_1[832967:829950]);
csa_3018 csau_3018_i138(A[1252469:1249452],A[1255487:1252470],A[1258505:1255488],tree_1[835985:832968],tree_1[839003:835986]);
csa_3018 csau_3018_i139(A[1261523:1258506],A[1264541:1261524],A[1267559:1264542],tree_1[842021:839004],tree_1[845039:842022]);
csa_3018 csau_3018_i140(A[1270577:1267560],A[1273595:1270578],A[1276613:1273596],tree_1[848057:845040],tree_1[851075:848058]);
csa_3018 csau_3018_i141(A[1279631:1276614],A[1282649:1279632],A[1285667:1282650],tree_1[854093:851076],tree_1[857111:854094]);
csa_3018 csau_3018_i142(A[1288685:1285668],A[1291703:1288686],A[1294721:1291704],tree_1[860129:857112],tree_1[863147:860130]);
csa_3018 csau_3018_i143(A[1297739:1294722],A[1300757:1297740],A[1303775:1300758],tree_1[866165:863148],tree_1[869183:866166]);
csa_3018 csau_3018_i144(A[1306793:1303776],A[1309811:1306794],A[1312829:1309812],tree_1[872201:869184],tree_1[875219:872202]);
csa_3018 csau_3018_i145(A[1315847:1312830],A[1318865:1315848],A[1321883:1318866],tree_1[878237:875220],tree_1[881255:878238]);
csa_3018 csau_3018_i146(A[1324901:1321884],A[1327919:1324902],A[1330937:1327920],tree_1[884273:881256],tree_1[887291:884274]);
csa_3018 csau_3018_i147(A[1333955:1330938],A[1336973:1333956],A[1339991:1336974],tree_1[890309:887292],tree_1[893327:890310]);
csa_3018 csau_3018_i148(A[1343009:1339992],A[1346027:1343010],A[1349045:1346028],tree_1[896345:893328],tree_1[899363:896346]);
csa_3018 csau_3018_i149(A[1352063:1349046],A[1355081:1352064],A[1358099:1355082],tree_1[902381:899364],tree_1[905399:902382]);
csa_3018 csau_3018_i150(A[1361117:1358100],A[1364135:1361118],A[1367153:1364136],tree_1[908417:905400],tree_1[911435:908418]);
csa_3018 csau_3018_i151(A[1370171:1367154],A[1373189:1370172],A[1376207:1373190],tree_1[914453:911436],tree_1[917471:914454]);
csa_3018 csau_3018_i152(A[1379225:1376208],A[1382243:1379226],A[1385261:1382244],tree_1[920489:917472],tree_1[923507:920490]);
csa_3018 csau_3018_i153(A[1388279:1385262],A[1391297:1388280],A[1394315:1391298],tree_1[926525:923508],tree_1[929543:926526]);
csa_3018 csau_3018_i154(A[1397333:1394316],A[1400351:1397334],A[1403369:1400352],tree_1[932561:929544],tree_1[935579:932562]);
csa_3018 csau_3018_i155(A[1406387:1403370],A[1409405:1406388],A[1412423:1409406],tree_1[938597:935580],tree_1[941615:938598]);
csa_3018 csau_3018_i156(A[1415441:1412424],A[1418459:1415442],A[1421477:1418460],tree_1[944633:941616],tree_1[947651:944634]);
csa_3018 csau_3018_i157(A[1424495:1421478],A[1427513:1424496],A[1430531:1427514],tree_1[950669:947652],tree_1[953687:950670]);
csa_3018 csau_3018_i158(A[1433549:1430532],A[1436567:1433550],A[1439585:1436568],tree_1[956705:953688],tree_1[959723:956706]);
csa_3018 csau_3018_i159(A[1442603:1439586],A[1445621:1442604],A[1448639:1445622],tree_1[962741:959724],tree_1[965759:962742]);
csa_3018 csau_3018_i160(A[1451657:1448640],A[1454675:1451658],A[1457693:1454676],tree_1[968777:965760],tree_1[971795:968778]);
csa_3018 csau_3018_i161(A[1460711:1457694],A[1463729:1460712],A[1466747:1463730],tree_1[974813:971796],tree_1[977831:974814]);
csa_3018 csau_3018_i162(A[1469765:1466748],A[1472783:1469766],A[1475801:1472784],tree_1[980849:977832],tree_1[983867:980850]);
csa_3018 csau_3018_i163(A[1478819:1475802],A[1481837:1478820],A[1484855:1481838],tree_1[986885:983868],tree_1[989903:986886]);
csa_3018 csau_3018_i164(A[1487873:1484856],A[1490891:1487874],A[1493909:1490892],tree_1[992921:989904],tree_1[995939:992922]);
csa_3018 csau_3018_i165(A[1496927:1493910],A[1499945:1496928],A[1502963:1499946],tree_1[998957:995940],tree_1[1001975:998958]);
csa_3018 csau_3018_i166(A[1505981:1502964],A[1508999:1505982],A[1512017:1509000],tree_1[1004993:1001976],tree_1[1008011:1004994]);
csa_3018 csau_3018_i167(A[1515035:1512018],A[1518053:1515036],A[1521071:1518054],tree_1[1011029:1008012],tree_1[1014047:1011030]);
csa_3018 csau_3018_i168(A[1524089:1521072],A[1527107:1524090],A[1530125:1527108],tree_1[1017065:1014048],tree_1[1020083:1017066]);
csa_3018 csau_3018_i169(A[1533143:1530126],A[1536161:1533144],A[1539179:1536162],tree_1[1023101:1020084],tree_1[1026119:1023102]);
csa_3018 csau_3018_i170(A[1542197:1539180],A[1545215:1542198],A[1548233:1545216],tree_1[1029137:1026120],tree_1[1032155:1029138]);
csa_3018 csau_3018_i171(A[1551251:1548234],A[1554269:1551252],A[1557287:1554270],tree_1[1035173:1032156],tree_1[1038191:1035174]);
csa_3018 csau_3018_i172(A[1560305:1557288],A[1563323:1560306],A[1566341:1563324],tree_1[1041209:1038192],tree_1[1044227:1041210]);
csa_3018 csau_3018_i173(A[1569359:1566342],A[1572377:1569360],A[1575395:1572378],tree_1[1047245:1044228],tree_1[1050263:1047246]);
csa_3018 csau_3018_i174(A[1578413:1575396],A[1581431:1578414],A[1584449:1581432],tree_1[1053281:1050264],tree_1[1056299:1053282]);
csa_3018 csau_3018_i175(A[1587467:1584450],A[1590485:1587468],A[1593503:1590486],tree_1[1059317:1056300],tree_1[1062335:1059318]);
csa_3018 csau_3018_i176(A[1596521:1593504],A[1599539:1596522],A[1602557:1599540],tree_1[1065353:1062336],tree_1[1068371:1065354]);
csa_3018 csau_3018_i177(A[1605575:1602558],A[1608593:1605576],A[1611611:1608594],tree_1[1071389:1068372],tree_1[1074407:1071390]);
csa_3018 csau_3018_i178(A[1614629:1611612],A[1617647:1614630],A[1620665:1617648],tree_1[1077425:1074408],tree_1[1080443:1077426]);
csa_3018 csau_3018_i179(A[1623683:1620666],A[1626701:1623684],A[1629719:1626702],tree_1[1083461:1080444],tree_1[1086479:1083462]);
csa_3018 csau_3018_i180(A[1632737:1629720],A[1635755:1632738],A[1638773:1635756],tree_1[1089497:1086480],tree_1[1092515:1089498]);
csa_3018 csau_3018_i181(A[1641791:1638774],A[1644809:1641792],A[1647827:1644810],tree_1[1095533:1092516],tree_1[1098551:1095534]);
csa_3018 csau_3018_i182(A[1650845:1647828],A[1653863:1650846],A[1656881:1653864],tree_1[1101569:1098552],tree_1[1104587:1101570]);
csa_3018 csau_3018_i183(A[1659899:1656882],A[1662917:1659900],A[1665935:1662918],tree_1[1107605:1104588],tree_1[1110623:1107606]);
csa_3018 csau_3018_i184(A[1668953:1665936],A[1671971:1668954],A[1674989:1671972],tree_1[1113641:1110624],tree_1[1116659:1113642]);
csa_3018 csau_3018_i185(A[1678007:1674990],A[1681025:1678008],A[1684043:1681026],tree_1[1119677:1116660],tree_1[1122695:1119678]);
csa_3018 csau_3018_i186(A[1687061:1684044],A[1690079:1687062],A[1693097:1690080],tree_1[1125713:1122696],tree_1[1128731:1125714]);
csa_3018 csau_3018_i187(A[1696115:1693098],A[1699133:1696116],A[1702151:1699134],tree_1[1131749:1128732],tree_1[1134767:1131750]);
csa_3018 csau_3018_i188(A[1705169:1702152],A[1708187:1705170],A[1711205:1708188],tree_1[1137785:1134768],tree_1[1140803:1137786]);
csa_3018 csau_3018_i189(A[1714223:1711206],A[1717241:1714224],A[1720259:1717242],tree_1[1143821:1140804],tree_1[1146839:1143822]);
csa_3018 csau_3018_i190(A[1723277:1720260],A[1726295:1723278],A[1729313:1726296],tree_1[1149857:1146840],tree_1[1152875:1149858]);
csa_3018 csau_3018_i191(A[1732331:1729314],A[1735349:1732332],A[1738367:1735350],tree_1[1155893:1152876],tree_1[1158911:1155894]);
csa_3018 csau_3018_i192(A[1741385:1738368],A[1744403:1741386],A[1747421:1744404],tree_1[1161929:1158912],tree_1[1164947:1161930]);
csa_3018 csau_3018_i193(A[1750439:1747422],A[1753457:1750440],A[1756475:1753458],tree_1[1167965:1164948],tree_1[1170983:1167966]);
csa_3018 csau_3018_i194(A[1759493:1756476],A[1762511:1759494],A[1765529:1762512],tree_1[1174001:1170984],tree_1[1177019:1174002]);
csa_3018 csau_3018_i195(A[1768547:1765530],A[1771565:1768548],A[1774583:1771566],tree_1[1180037:1177020],tree_1[1183055:1180038]);
csa_3018 csau_3018_i196(A[1777601:1774584],A[1780619:1777602],A[1783637:1780620],tree_1[1186073:1183056],tree_1[1189091:1186074]);
csa_3018 csau_3018_i197(A[1786655:1783638],A[1789673:1786656],A[1792691:1789674],tree_1[1192109:1189092],tree_1[1195127:1192110]);
csa_3018 csau_3018_i198(A[1795709:1792692],A[1798727:1795710],A[1801745:1798728],tree_1[1198145:1195128],tree_1[1201163:1198146]);
csa_3018 csau_3018_i199(A[1804763:1801746],A[1807781:1804764],A[1810799:1807782],tree_1[1204181:1201164],tree_1[1207199:1204182]);
csa_3018 csau_3018_i200(A[1813817:1810800],A[1816835:1813818],A[1819853:1816836],tree_1[1210217:1207200],tree_1[1213235:1210218]);
csa_3018 csau_3018_i201(A[1822871:1819854],A[1825889:1822872],A[1828907:1825890],tree_1[1216253:1213236],tree_1[1219271:1216254]);
csa_3018 csau_3018_i202(A[1831925:1828908],A[1834943:1831926],A[1837961:1834944],tree_1[1222289:1219272],tree_1[1225307:1222290]);
csa_3018 csau_3018_i203(A[1840979:1837962],A[1843997:1840980],A[1847015:1843998],tree_1[1228325:1225308],tree_1[1231343:1228326]);
csa_3018 csau_3018_i204(A[1850033:1847016],A[1853051:1850034],A[1856069:1853052],tree_1[1234361:1231344],tree_1[1237379:1234362]);
csa_3018 csau_3018_i205(A[1859087:1856070],A[1862105:1859088],A[1865123:1862106],tree_1[1240397:1237380],tree_1[1243415:1240398]);
csa_3018 csau_3018_i206(A[1868141:1865124],A[1871159:1868142],A[1874177:1871160],tree_1[1246433:1243416],tree_1[1249451:1246434]);
csa_3018 csau_3018_i207(A[1877195:1874178],A[1880213:1877196],A[1883231:1880214],tree_1[1252469:1249452],tree_1[1255487:1252470]);
csa_3018 csau_3018_i208(A[1886249:1883232],A[1889267:1886250],A[1892285:1889268],tree_1[1258505:1255488],tree_1[1261523:1258506]);
csa_3018 csau_3018_i209(A[1895303:1892286],A[1898321:1895304],A[1901339:1898322],tree_1[1264541:1261524],tree_1[1267559:1264542]);
csa_3018 csau_3018_i210(A[1904357:1901340],A[1907375:1904358],A[1910393:1907376],tree_1[1270577:1267560],tree_1[1273595:1270578]);
csa_3018 csau_3018_i211(A[1913411:1910394],A[1916429:1913412],A[1919447:1916430],tree_1[1276613:1273596],tree_1[1279631:1276614]);
csa_3018 csau_3018_i212(A[1922465:1919448],A[1925483:1922466],A[1928501:1925484],tree_1[1282649:1279632],tree_1[1285667:1282650]);
csa_3018 csau_3018_i213(A[1931519:1928502],A[1934537:1931520],A[1937555:1934538],tree_1[1288685:1285668],tree_1[1291703:1288686]);
csa_3018 csau_3018_i214(A[1940573:1937556],A[1943591:1940574],A[1946609:1943592],tree_1[1294721:1291704],tree_1[1297739:1294722]);
csa_3018 csau_3018_i215(A[1949627:1946610],A[1952645:1949628],A[1955663:1952646],tree_1[1300757:1297740],tree_1[1303775:1300758]);
csa_3018 csau_3018_i216(A[1958681:1955664],A[1961699:1958682],A[1964717:1961700],tree_1[1306793:1303776],tree_1[1309811:1306794]);
csa_3018 csau_3018_i217(A[1967735:1964718],A[1970753:1967736],A[1973771:1970754],tree_1[1312829:1309812],tree_1[1315847:1312830]);
csa_3018 csau_3018_i218(A[1976789:1973772],A[1979807:1976790],A[1982825:1979808],tree_1[1318865:1315848],tree_1[1321883:1318866]);
csa_3018 csau_3018_i219(A[1985843:1982826],A[1988861:1985844],A[1991879:1988862],tree_1[1324901:1321884],tree_1[1327919:1324902]);
csa_3018 csau_3018_i220(A[1994897:1991880],A[1997915:1994898],A[2000933:1997916],tree_1[1330937:1327920],tree_1[1333955:1330938]);
csa_3018 csau_3018_i221(A[2003951:2000934],A[2006969:2003952],A[2009987:2006970],tree_1[1336973:1333956],tree_1[1339991:1336974]);
csa_3018 csau_3018_i222(A[2013005:2009988],A[2016023:2013006],A[2019041:2016024],tree_1[1343009:1339992],tree_1[1346027:1343010]);
csa_3018 csau_3018_i223(A[2022059:2019042],A[2025077:2022060],A[2028095:2025078],tree_1[1349045:1346028],tree_1[1352063:1349046]);
csa_3018 csau_3018_i224(A[2031113:2028096],A[2034131:2031114],A[2037149:2034132],tree_1[1355081:1352064],tree_1[1358099:1355082]);
csa_3018 csau_3018_i225(A[2040167:2037150],A[2043185:2040168],A[2046203:2043186],tree_1[1361117:1358100],tree_1[1364135:1361118]);
csa_3018 csau_3018_i226(A[2049221:2046204],A[2052239:2049222],A[2055257:2052240],tree_1[1367153:1364136],tree_1[1370171:1367154]);
csa_3018 csau_3018_i227(A[2058275:2055258],A[2061293:2058276],A[2064311:2061294],tree_1[1373189:1370172],tree_1[1376207:1373190]);
csa_3018 csau_3018_i228(A[2067329:2064312],A[2070347:2067330],A[2073365:2070348],tree_1[1379225:1376208],tree_1[1382243:1379226]);
csa_3018 csau_3018_i229(A[2076383:2073366],A[2079401:2076384],A[2082419:2079402],tree_1[1385261:1382244],tree_1[1388279:1385262]);
csa_3018 csau_3018_i230(A[2085437:2082420],A[2088455:2085438],A[2091473:2088456],tree_1[1391297:1388280],tree_1[1394315:1391298]);
csa_3018 csau_3018_i231(A[2094491:2091474],A[2097509:2094492],A[2100527:2097510],tree_1[1397333:1394316],tree_1[1400351:1397334]);
csa_3018 csau_3018_i232(A[2103545:2100528],A[2106563:2103546],A[2109581:2106564],tree_1[1403369:1400352],tree_1[1406387:1403370]);
csa_3018 csau_3018_i233(A[2112599:2109582],A[2115617:2112600],A[2118635:2115618],tree_1[1409405:1406388],tree_1[1412423:1409406]);
csa_3018 csau_3018_i234(A[2121653:2118636],A[2124671:2121654],A[2127689:2124672],tree_1[1415441:1412424],tree_1[1418459:1415442]);
csa_3018 csau_3018_i235(A[2130707:2127690],A[2133725:2130708],A[2136743:2133726],tree_1[1421477:1418460],tree_1[1424495:1421478]);
csa_3018 csau_3018_i236(A[2139761:2136744],A[2142779:2139762],A[2145797:2142780],tree_1[1427513:1424496],tree_1[1430531:1427514]);
csa_3018 csau_3018_i237(A[2148815:2145798],A[2151833:2148816],A[2154851:2151834],tree_1[1433549:1430532],tree_1[1436567:1433550]);
csa_3018 csau_3018_i238(A[2157869:2154852],A[2160887:2157870],A[2163905:2160888],tree_1[1439585:1436568],tree_1[1442603:1439586]);
csa_3018 csau_3018_i239(A[2166923:2163906],A[2169941:2166924],A[2172959:2169942],tree_1[1445621:1442604],tree_1[1448639:1445622]);
csa_3018 csau_3018_i240(A[2175977:2172960],A[2178995:2175978],A[2182013:2178996],tree_1[1451657:1448640],tree_1[1454675:1451658]);
csa_3018 csau_3018_i241(A[2185031:2182014],A[2188049:2185032],A[2191067:2188050],tree_1[1457693:1454676],tree_1[1460711:1457694]);
csa_3018 csau_3018_i242(A[2194085:2191068],A[2197103:2194086],A[2200121:2197104],tree_1[1463729:1460712],tree_1[1466747:1463730]);
csa_3018 csau_3018_i243(A[2203139:2200122],A[2206157:2203140],A[2209175:2206158],tree_1[1469765:1466748],tree_1[1472783:1469766]);
csa_3018 csau_3018_i244(A[2212193:2209176],A[2215211:2212194],A[2218229:2215212],tree_1[1475801:1472784],tree_1[1478819:1475802]);
csa_3018 csau_3018_i245(A[2221247:2218230],A[2224265:2221248],A[2227283:2224266],tree_1[1481837:1478820],tree_1[1484855:1481838]);
csa_3018 csau_3018_i246(A[2230301:2227284],A[2233319:2230302],A[2236337:2233320],tree_1[1487873:1484856],tree_1[1490891:1487874]);
csa_3018 csau_3018_i247(A[2239355:2236338],A[2242373:2239356],A[2245391:2242374],tree_1[1493909:1490892],tree_1[1496927:1493910]);
csa_3018 csau_3018_i248(A[2248409:2245392],A[2251427:2248410],A[2254445:2251428],tree_1[1499945:1496928],tree_1[1502963:1499946]);
csa_3018 csau_3018_i249(A[2257463:2254446],A[2260481:2257464],A[2263499:2260482],tree_1[1505981:1502964],tree_1[1508999:1505982]);
csa_3018 csau_3018_i250(A[2266517:2263500],A[2269535:2266518],A[2272553:2269536],tree_1[1512017:1509000],tree_1[1515035:1512018]);
csa_3018 csau_3018_i251(A[2275571:2272554],A[2278589:2275572],A[2281607:2278590],tree_1[1518053:1515036],tree_1[1521071:1518054]);
csa_3018 csau_3018_i252(A[2284625:2281608],A[2287643:2284626],A[2290661:2287644],tree_1[1524089:1521072],tree_1[1527107:1524090]);
csa_3018 csau_3018_i253(A[2293679:2290662],A[2296697:2293680],A[2299715:2296698],tree_1[1530125:1527108],tree_1[1533143:1530126]);
csa_3018 csau_3018_i254(A[2302733:2299716],A[2305751:2302734],A[2308769:2305752],tree_1[1536161:1533144],tree_1[1539179:1536162]);
csa_3018 csau_3018_i255(A[2311787:2308770],A[2314805:2311788],A[2317823:2314806],tree_1[1542197:1539180],tree_1[1545215:1542198]);
csa_3018 csau_3018_i256(A[2320841:2317824],A[2323859:2320842],A[2326877:2323860],tree_1[1548233:1545216],tree_1[1551251:1548234]);
csa_3018 csau_3018_i257(A[2329895:2326878],A[2332913:2329896],A[2335931:2332914],tree_1[1554269:1551252],tree_1[1557287:1554270]);
csa_3018 csau_3018_i258(A[2338949:2335932],A[2341967:2338950],A[2344985:2341968],tree_1[1560305:1557288],tree_1[1563323:1560306]);
csa_3018 csau_3018_i259(A[2348003:2344986],A[2351021:2348004],A[2354039:2351022],tree_1[1566341:1563324],tree_1[1569359:1566342]);
csa_3018 csau_3018_i260(A[2357057:2354040],A[2360075:2357058],A[2363093:2360076],tree_1[1572377:1569360],tree_1[1575395:1572378]);
csa_3018 csau_3018_i261(A[2366111:2363094],A[2369129:2366112],A[2372147:2369130],tree_1[1578413:1575396],tree_1[1581431:1578414]);
csa_3018 csau_3018_i262(A[2375165:2372148],A[2378183:2375166],A[2381201:2378184],tree_1[1584449:1581432],tree_1[1587467:1584450]);
csa_3018 csau_3018_i263(A[2384219:2381202],A[2387237:2384220],A[2390255:2387238],tree_1[1590485:1587468],tree_1[1593503:1590486]);
csa_3018 csau_3018_i264(A[2393273:2390256],A[2396291:2393274],A[2399309:2396292],tree_1[1596521:1593504],tree_1[1599539:1596522]);
csa_3018 csau_3018_i265(A[2402327:2399310],A[2405345:2402328],A[2408363:2405346],tree_1[1602557:1599540],tree_1[1605575:1602558]);
csa_3018 csau_3018_i266(A[2411381:2408364],A[2414399:2411382],A[2417417:2414400],tree_1[1608593:1605576],tree_1[1611611:1608594]);
csa_3018 csau_3018_i267(A[2420435:2417418],A[2423453:2420436],A[2426471:2423454],tree_1[1614629:1611612],tree_1[1617647:1614630]);
csa_3018 csau_3018_i268(A[2429489:2426472],A[2432507:2429490],A[2435525:2432508],tree_1[1620665:1617648],tree_1[1623683:1620666]);
csa_3018 csau_3018_i269(A[2438543:2435526],A[2441561:2438544],A[2444579:2441562],tree_1[1626701:1623684],tree_1[1629719:1626702]);
csa_3018 csau_3018_i270(A[2447597:2444580],A[2450615:2447598],A[2453633:2450616],tree_1[1632737:1629720],tree_1[1635755:1632738]);
csa_3018 csau_3018_i271(A[2456651:2453634],A[2459669:2456652],A[2462687:2459670],tree_1[1638773:1635756],tree_1[1641791:1638774]);
csa_3018 csau_3018_i272(A[2465705:2462688],A[2468723:2465706],A[2471741:2468724],tree_1[1644809:1641792],tree_1[1647827:1644810]);
csa_3018 csau_3018_i273(A[2474759:2471742],A[2477777:2474760],A[2480795:2477778],tree_1[1650845:1647828],tree_1[1653863:1650846]);
csa_3018 csau_3018_i274(A[2483813:2480796],A[2486831:2483814],A[2489849:2486832],tree_1[1656881:1653864],tree_1[1659899:1656882]);
csa_3018 csau_3018_i275(A[2492867:2489850],A[2495885:2492868],A[2498903:2495886],tree_1[1662917:1659900],tree_1[1665935:1662918]);
csa_3018 csau_3018_i276(A[2501921:2498904],A[2504939:2501922],A[2507957:2504940],tree_1[1668953:1665936],tree_1[1671971:1668954]);
csa_3018 csau_3018_i277(A[2510975:2507958],A[2513993:2510976],A[2517011:2513994],tree_1[1674989:1671972],tree_1[1678007:1674990]);
csa_3018 csau_3018_i278(A[2520029:2517012],A[2523047:2520030],A[2526065:2523048],tree_1[1681025:1678008],tree_1[1684043:1681026]);
csa_3018 csau_3018_i279(A[2529083:2526066],A[2532101:2529084],A[2535119:2532102],tree_1[1687061:1684044],tree_1[1690079:1687062]);
csa_3018 csau_3018_i280(A[2538137:2535120],A[2541155:2538138],A[2544173:2541156],tree_1[1693097:1690080],tree_1[1696115:1693098]);
csa_3018 csau_3018_i281(A[2547191:2544174],A[2550209:2547192],A[2553227:2550210],tree_1[1699133:1696116],tree_1[1702151:1699134]);
csa_3018 csau_3018_i282(A[2556245:2553228],A[2559263:2556246],A[2562281:2559264],tree_1[1705169:1702152],tree_1[1708187:1705170]);
csa_3018 csau_3018_i283(A[2565299:2562282],A[2568317:2565300],A[2571335:2568318],tree_1[1711205:1708188],tree_1[1714223:1711206]);
csa_3018 csau_3018_i284(A[2574353:2571336],A[2577371:2574354],A[2580389:2577372],tree_1[1717241:1714224],tree_1[1720259:1717242]);
csa_3018 csau_3018_i285(A[2583407:2580390],A[2586425:2583408],A[2589443:2586426],tree_1[1723277:1720260],tree_1[1726295:1723278]);
csa_3018 csau_3018_i286(A[2592461:2589444],A[2595479:2592462],A[2598497:2595480],tree_1[1729313:1726296],tree_1[1732331:1729314]);
csa_3018 csau_3018_i287(A[2601515:2598498],A[2604533:2601516],A[2607551:2604534],tree_1[1735349:1732332],tree_1[1738367:1735350]);
csa_3018 csau_3018_i288(A[2610569:2607552],A[2613587:2610570],A[2616605:2613588],tree_1[1741385:1738368],tree_1[1744403:1741386]);
csa_3018 csau_3018_i289(A[2619623:2616606],A[2622641:2619624],A[2625659:2622642],tree_1[1747421:1744404],tree_1[1750439:1747422]);
csa_3018 csau_3018_i290(A[2628677:2625660],A[2631695:2628678],A[2634713:2631696],tree_1[1753457:1750440],tree_1[1756475:1753458]);
csa_3018 csau_3018_i291(A[2637731:2634714],A[2640749:2637732],A[2643767:2640750],tree_1[1759493:1756476],tree_1[1762511:1759494]);
csa_3018 csau_3018_i292(A[2646785:2643768],A[2649803:2646786],A[2652821:2649804],tree_1[1765529:1762512],tree_1[1768547:1765530]);
csa_3018 csau_3018_i293(A[2655839:2652822],A[2658857:2655840],A[2661875:2658858],tree_1[1771565:1768548],tree_1[1774583:1771566]);
csa_3018 csau_3018_i294(A[2664893:2661876],A[2667911:2664894],A[2670929:2667912],tree_1[1777601:1774584],tree_1[1780619:1777602]);
csa_3018 csau_3018_i295(A[2673947:2670930],A[2676965:2673948],A[2679983:2676966],tree_1[1783637:1780620],tree_1[1786655:1783638]);
csa_3018 csau_3018_i296(A[2683001:2679984],A[2686019:2683002],A[2689037:2686020],tree_1[1789673:1786656],tree_1[1792691:1789674]);
csa_3018 csau_3018_i297(A[2692055:2689038],A[2695073:2692056],A[2698091:2695074],tree_1[1795709:1792692],tree_1[1798727:1795710]);
csa_3018 csau_3018_i298(A[2701109:2698092],A[2704127:2701110],A[2707145:2704128],tree_1[1801745:1798728],tree_1[1804763:1801746]);
csa_3018 csau_3018_i299(A[2710163:2707146],A[2713181:2710164],A[2716199:2713182],tree_1[1807781:1804764],tree_1[1810799:1807782]);
csa_3018 csau_3018_i300(A[2719217:2716200],A[2722235:2719218],A[2725253:2722236],tree_1[1813817:1810800],tree_1[1816835:1813818]);
csa_3018 csau_3018_i301(A[2728271:2725254],A[2731289:2728272],A[2734307:2731290],tree_1[1819853:1816836],tree_1[1822871:1819854]);
csa_3018 csau_3018_i302(A[2737325:2734308],A[2740343:2737326],A[2743361:2740344],tree_1[1825889:1822872],tree_1[1828907:1825890]);
csa_3018 csau_3018_i303(A[2746379:2743362],A[2749397:2746380],A[2752415:2749398],tree_1[1831925:1828908],tree_1[1834943:1831926]);
csa_3018 csau_3018_i304(A[2755433:2752416],A[2758451:2755434],A[2761469:2758452],tree_1[1837961:1834944],tree_1[1840979:1837962]);
csa_3018 csau_3018_i305(A[2764487:2761470],A[2767505:2764488],A[2770523:2767506],tree_1[1843997:1840980],tree_1[1847015:1843998]);
csa_3018 csau_3018_i306(A[2773541:2770524],A[2776559:2773542],A[2779577:2776560],tree_1[1850033:1847016],tree_1[1853051:1850034]);
csa_3018 csau_3018_i307(A[2782595:2779578],A[2785613:2782596],A[2788631:2785614],tree_1[1856069:1853052],tree_1[1859087:1856070]);
csa_3018 csau_3018_i308(A[2791649:2788632],A[2794667:2791650],A[2797685:2794668],tree_1[1862105:1859088],tree_1[1865123:1862106]);
csa_3018 csau_3018_i309(A[2800703:2797686],A[2803721:2800704],A[2806739:2803722],tree_1[1868141:1865124],tree_1[1871159:1868142]);
csa_3018 csau_3018_i310(A[2809757:2806740],A[2812775:2809758],A[2815793:2812776],tree_1[1874177:1871160],tree_1[1877195:1874178]);
csa_3018 csau_3018_i311(A[2818811:2815794],A[2821829:2818812],A[2824847:2821830],tree_1[1880213:1877196],tree_1[1883231:1880214]);
csa_3018 csau_3018_i312(A[2827865:2824848],A[2830883:2827866],A[2833901:2830884],tree_1[1886249:1883232],tree_1[1889267:1886250]);
csa_3018 csau_3018_i313(A[2836919:2833902],A[2839937:2836920],A[2842955:2839938],tree_1[1892285:1889268],tree_1[1895303:1892286]);
csa_3018 csau_3018_i314(A[2845973:2842956],A[2848991:2845974],A[2852009:2848992],tree_1[1898321:1895304],tree_1[1901339:1898322]);
csa_3018 csau_3018_i315(A[2855027:2852010],A[2858045:2855028],A[2861063:2858046],tree_1[1904357:1901340],tree_1[1907375:1904358]);
csa_3018 csau_3018_i316(A[2864081:2861064],A[2867099:2864082],A[2870117:2867100],tree_1[1910393:1907376],tree_1[1913411:1910394]);
csa_3018 csau_3018_i317(A[2873135:2870118],A[2876153:2873136],A[2879171:2876154],tree_1[1916429:1913412],tree_1[1919447:1916430]);
csa_3018 csau_3018_i318(A[2882189:2879172],A[2885207:2882190],A[2888225:2885208],tree_1[1922465:1919448],tree_1[1925483:1922466]);
csa_3018 csau_3018_i319(A[2891243:2888226],A[2894261:2891244],A[2897279:2894262],tree_1[1928501:1925484],tree_1[1931519:1928502]);
csa_3018 csau_3018_i320(A[2900297:2897280],A[2903315:2900298],A[2906333:2903316],tree_1[1934537:1931520],tree_1[1937555:1934538]);
csa_3018 csau_3018_i321(A[2909351:2906334],A[2912369:2909352],A[2915387:2912370],tree_1[1940573:1937556],tree_1[1943591:1940574]);
csa_3018 csau_3018_i322(A[2918405:2915388],A[2921423:2918406],A[2924441:2921424],tree_1[1946609:1943592],tree_1[1949627:1946610]);
csa_3018 csau_3018_i323(A[2927459:2924442],A[2930477:2927460],A[2933495:2930478],tree_1[1952645:1949628],tree_1[1955663:1952646]);
csa_3018 csau_3018_i324(A[2936513:2933496],A[2939531:2936514],A[2942549:2939532],tree_1[1958681:1955664],tree_1[1961699:1958682]);
csa_3018 csau_3018_i325(A[2945567:2942550],A[2948585:2945568],A[2951603:2948586],tree_1[1964717:1961700],tree_1[1967735:1964718]);
csa_3018 csau_3018_i326(A[2954621:2951604],A[2957639:2954622],A[2960657:2957640],tree_1[1970753:1967736],tree_1[1973771:1970754]);
csa_3018 csau_3018_i327(A[2963675:2960658],A[2966693:2963676],A[2969711:2966694],tree_1[1976789:1973772],tree_1[1979807:1976790]);
csa_3018 csau_3018_i328(A[2972729:2969712],A[2975747:2972730],A[2978765:2975748],tree_1[1982825:1979808],tree_1[1985843:1982826]);
csa_3018 csau_3018_i329(A[2981783:2978766],A[2984801:2981784],A[2987819:2984802],tree_1[1988861:1985844],tree_1[1991879:1988862]);
csa_3018 csau_3018_i330(A[2990837:2987820],A[2993855:2990838],A[2996873:2993856],tree_1[1994897:1991880],tree_1[1997915:1994898]);
csa_3018 csau_3018_i331(A[2999891:2996874],A[3002909:2999892],A[3005927:3002910],tree_1[2000933:1997916],tree_1[2003951:2000934]);
csa_3018 csau_3018_i332(A[3008945:3005928],A[3011963:3008946],A[3014981:3011964],tree_1[2006969:2003952],tree_1[2009987:2006970]);
csa_3018 csau_3018_i333(A[3017999:3014982],A[3021017:3018000],A[3024035:3021018],tree_1[2013005:2009988],tree_1[2016023:2013006]);
csa_3018 csau_3018_i334(A[3027053:3024036],A[3030071:3027054],A[3033089:3030072],tree_1[2019041:2016024],tree_1[2022059:2019042]);
csa_3018 csau_3018_i335(A[3036107:3033090],A[3039125:3036108],A[3042143:3039126],tree_1[2025077:2022060],tree_1[2028095:2025078]);
csa_3018 csau_3018_i336(A[3045161:3042144],A[3048179:3045162],A[3051197:3048180],tree_1[2031113:2028096],tree_1[2034131:2031114]);
csa_3018 csau_3018_i337(A[3054215:3051198],A[3057233:3054216],A[3060251:3057234],tree_1[2037149:2034132],tree_1[2040167:2037150]);
csa_3018 csau_3018_i338(A[3063269:3060252],A[3066287:3063270],A[3069305:3066288],tree_1[2043185:2040168],tree_1[2046203:2043186]);
csa_3018 csau_3018_i339(A[3072323:3069306],A[3075341:3072324],A[3078359:3075342],tree_1[2049221:2046204],tree_1[2052239:2049222]);
csa_3018 csau_3018_i340(A[3081377:3078360],A[3084395:3081378],A[3087413:3084396],tree_1[2055257:2052240],tree_1[2058275:2055258]);
csa_3018 csau_3018_i341(A[3090431:3087414],A[3093449:3090432],A[3096467:3093450],tree_1[2061293:2058276],tree_1[2064311:2061294]);
csa_3018 csau_3018_i342(A[3099485:3096468],A[3102503:3099486],A[3105521:3102504],tree_1[2067329:2064312],tree_1[2070347:2067330]);
csa_3018 csau_3018_i343(A[3108539:3105522],A[3111557:3108540],A[3114575:3111558],tree_1[2073365:2070348],tree_1[2076383:2073366]);
csa_3018 csau_3018_i344(A[3117593:3114576],A[3120611:3117594],A[3123629:3120612],tree_1[2079401:2076384],tree_1[2082419:2079402]);
csa_3018 csau_3018_i345(A[3126647:3123630],A[3129665:3126648],A[3132683:3129666],tree_1[2085437:2082420],tree_1[2088455:2085438]);
csa_3018 csau_3018_i346(A[3135701:3132684],A[3138719:3135702],A[3141737:3138720],tree_1[2091473:2088456],tree_1[2094491:2091474]);
csa_3018 csau_3018_i347(A[3144755:3141738],A[3147773:3144756],A[3150791:3147774],tree_1[2097509:2094492],tree_1[2100527:2097510]);
csa_3018 csau_3018_i348(A[3153809:3150792],A[3156827:3153810],A[3159845:3156828],tree_1[2103545:2100528],tree_1[2106563:2103546]);
csa_3018 csau_3018_i349(A[3162863:3159846],A[3165881:3162864],A[3168899:3165882],tree_1[2109581:2106564],tree_1[2112599:2109582]);
csa_3018 csau_3018_i350(A[3171917:3168900],A[3174935:3171918],A[3177953:3174936],tree_1[2115617:2112600],tree_1[2118635:2115618]);
csa_3018 csau_3018_i351(A[3180971:3177954],A[3183989:3180972],A[3187007:3183990],tree_1[2121653:2118636],tree_1[2124671:2121654]);
csa_3018 csau_3018_i352(A[3190025:3187008],A[3193043:3190026],A[3196061:3193044],tree_1[2127689:2124672],tree_1[2130707:2127690]);
csa_3018 csau_3018_i353(A[3199079:3196062],A[3202097:3199080],A[3205115:3202098],tree_1[2133725:2130708],tree_1[2136743:2133726]);
csa_3018 csau_3018_i354(A[3208133:3205116],A[3211151:3208134],A[3214169:3211152],tree_1[2139761:2136744],tree_1[2142779:2139762]);
csa_3018 csau_3018_i355(A[3217187:3214170],A[3220205:3217188],A[3223223:3220206],tree_1[2145797:2142780],tree_1[2148815:2145798]);
csa_3018 csau_3018_i356(A[3226241:3223224],A[3229259:3226242],A[3232277:3229260],tree_1[2151833:2148816],tree_1[2154851:2151834]);
csa_3018 csau_3018_i357(A[3235295:3232278],A[3238313:3235296],A[3241331:3238314],tree_1[2157869:2154852],tree_1[2160887:2157870]);
csa_3018 csau_3018_i358(A[3244349:3241332],A[3247367:3244350],A[3250385:3247368],tree_1[2163905:2160888],tree_1[2166923:2163906]);
csa_3018 csau_3018_i359(A[3253403:3250386],A[3256421:3253404],A[3259439:3256422],tree_1[2169941:2166924],tree_1[2172959:2169942]);
csa_3018 csau_3018_i360(A[3262457:3259440],A[3265475:3262458],A[3268493:3265476],tree_1[2175977:2172960],tree_1[2178995:2175978]);
csa_3018 csau_3018_i361(A[3271511:3268494],A[3274529:3271512],A[3277547:3274530],tree_1[2182013:2178996],tree_1[2185031:2182014]);
csa_3018 csau_3018_i362(A[3280565:3277548],A[3283583:3280566],A[3286601:3283584],tree_1[2188049:2185032],tree_1[2191067:2188050]);
csa_3018 csau_3018_i363(A[3289619:3286602],A[3292637:3289620],A[3295655:3292638],tree_1[2194085:2191068],tree_1[2197103:2194086]);
csa_3018 csau_3018_i364(A[3298673:3295656],A[3301691:3298674],A[3304709:3301692],tree_1[2200121:2197104],tree_1[2203139:2200122]);
csa_3018 csau_3018_i365(A[3307727:3304710],A[3310745:3307728],A[3313763:3310746],tree_1[2206157:2203140],tree_1[2209175:2206158]);
csa_3018 csau_3018_i366(A[3316781:3313764],A[3319799:3316782],A[3322817:3319800],tree_1[2212193:2209176],tree_1[2215211:2212194]);
csa_3018 csau_3018_i367(A[3325835:3322818],A[3328853:3325836],A[3331871:3328854],tree_1[2218229:2215212],tree_1[2221247:2218230]);
csa_3018 csau_3018_i368(A[3334889:3331872],A[3337907:3334890],A[3340925:3337908],tree_1[2224265:2221248],tree_1[2227283:2224266]);
csa_3018 csau_3018_i369(A[3343943:3340926],A[3346961:3343944],A[3349979:3346962],tree_1[2230301:2227284],tree_1[2233319:2230302]);
csa_3018 csau_3018_i370(A[3352997:3349980],A[3356015:3352998],A[3359033:3356016],tree_1[2236337:2233320],tree_1[2239355:2236338]);
csa_3018 csau_3018_i371(A[3362051:3359034],A[3365069:3362052],A[3368087:3365070],tree_1[2242373:2239356],tree_1[2245391:2242374]);
csa_3018 csau_3018_i372(A[3371105:3368088],A[3374123:3371106],A[3377141:3374124],tree_1[2248409:2245392],tree_1[2251427:2248410]);
csa_3018 csau_3018_i373(A[3380159:3377142],A[3383177:3380160],A[3386195:3383178],tree_1[2254445:2251428],tree_1[2257463:2254446]);
csa_3018 csau_3018_i374(A[3389213:3386196],A[3392231:3389214],A[3395249:3392232],tree_1[2260481:2257464],tree_1[2263499:2260482]);
csa_3018 csau_3018_i375(A[3398267:3395250],A[3401285:3398268],A[3404303:3401286],tree_1[2266517:2263500],tree_1[2269535:2266518]);
csa_3018 csau_3018_i376(A[3407321:3404304],A[3410339:3407322],A[3413357:3410340],tree_1[2272553:2269536],tree_1[2275571:2272554]);
csa_3018 csau_3018_i377(A[3416375:3413358],A[3419393:3416376],A[3422411:3419394],tree_1[2278589:2275572],tree_1[2281607:2278590]);
csa_3018 csau_3018_i378(A[3425429:3422412],A[3428447:3425430],A[3431465:3428448],tree_1[2284625:2281608],tree_1[2287643:2284626]);
csa_3018 csau_3018_i379(A[3434483:3431466],A[3437501:3434484],A[3440519:3437502],tree_1[2290661:2287644],tree_1[2293679:2290662]);
csa_3018 csau_3018_i380(A[3443537:3440520],A[3446555:3443538],A[3449573:3446556],tree_1[2296697:2293680],tree_1[2299715:2296698]);
csa_3018 csau_3018_i381(A[3452591:3449574],A[3455609:3452592],A[3458627:3455610],tree_1[2302733:2299716],tree_1[2305751:2302734]);
csa_3018 csau_3018_i382(A[3461645:3458628],A[3464663:3461646],A[3467681:3464664],tree_1[2308769:2305752],tree_1[2311787:2308770]);
csa_3018 csau_3018_i383(A[3470699:3467682],A[3473717:3470700],A[3476735:3473718],tree_1[2314805:2311788],tree_1[2317823:2314806]);
csa_3018 csau_3018_i384(A[3479753:3476736],A[3482771:3479754],A[3485789:3482772],tree_1[2320841:2317824],tree_1[2323859:2320842]);
csa_3018 csau_3018_i385(A[3488807:3485790],A[3491825:3488808],A[3494843:3491826],tree_1[2326877:2323860],tree_1[2329895:2326878]);
csa_3018 csau_3018_i386(A[3497861:3494844],A[3500879:3497862],A[3503897:3500880],tree_1[2332913:2329896],tree_1[2335931:2332914]);
csa_3018 csau_3018_i387(A[3506915:3503898],A[3509933:3506916],A[3512951:3509934],tree_1[2338949:2335932],tree_1[2341967:2338950]);
csa_3018 csau_3018_i388(A[3515969:3512952],A[3518987:3515970],A[3522005:3518988],tree_1[2344985:2341968],tree_1[2348003:2344986]);
csa_3018 csau_3018_i389(A[3525023:3522006],A[3528041:3525024],A[3531059:3528042],tree_1[2351021:2348004],tree_1[2354039:2351022]);
csa_3018 csau_3018_i390(A[3534077:3531060],A[3537095:3534078],A[3540113:3537096],tree_1[2357057:2354040],tree_1[2360075:2357058]);
csa_3018 csau_3018_i391(A[3543131:3540114],A[3546149:3543132],A[3549167:3546150],tree_1[2363093:2360076],tree_1[2366111:2363094]);
csa_3018 csau_3018_i392(A[3552185:3549168],A[3555203:3552186],A[3558221:3555204],tree_1[2369129:2366112],tree_1[2372147:2369130]);
csa_3018 csau_3018_i393(A[3561239:3558222],A[3564257:3561240],A[3567275:3564258],tree_1[2375165:2372148],tree_1[2378183:2375166]);
csa_3018 csau_3018_i394(A[3570293:3567276],A[3573311:3570294],A[3576329:3573312],tree_1[2381201:2378184],tree_1[2384219:2381202]);
csa_3018 csau_3018_i395(A[3579347:3576330],A[3582365:3579348],A[3585383:3582366],tree_1[2387237:2384220],tree_1[2390255:2387238]);
csa_3018 csau_3018_i396(A[3588401:3585384],A[3591419:3588402],A[3594437:3591420],tree_1[2393273:2390256],tree_1[2396291:2393274]);
csa_3018 csau_3018_i397(A[3597455:3594438],A[3600473:3597456],A[3603491:3600474],tree_1[2399309:2396292],tree_1[2402327:2399310]);
csa_3018 csau_3018_i398(A[3606509:3603492],A[3609527:3606510],A[3612545:3609528],tree_1[2405345:2402328],tree_1[2408363:2405346]);
csa_3018 csau_3018_i399(A[3615563:3612546],A[3618581:3615564],A[3621599:3618582],tree_1[2411381:2408364],tree_1[2414399:2411382]);
csa_3018 csau_3018_i400(A[3624617:3621600],A[3627635:3624618],A[3630653:3627636],tree_1[2417417:2414400],tree_1[2420435:2417418]);
csa_3018 csau_3018_i401(A[3633671:3630654],A[3636689:3633672],A[3639707:3636690],tree_1[2423453:2420436],tree_1[2426471:2423454]);
csa_3018 csau_3018_i402(A[3642725:3639708],A[3645743:3642726],A[3648761:3645744],tree_1[2429489:2426472],tree_1[2432507:2429490]);
csa_3018 csau_3018_i403(A[3651779:3648762],A[3654797:3651780],A[3657815:3654798],tree_1[2435525:2432508],tree_1[2438543:2435526]);
csa_3018 csau_3018_i404(A[3660833:3657816],A[3663851:3660834],A[3666869:3663852],tree_1[2441561:2438544],tree_1[2444579:2441562]);
csa_3018 csau_3018_i405(A[3669887:3666870],A[3672905:3669888],A[3675923:3672906],tree_1[2447597:2444580],tree_1[2450615:2447598]);
csa_3018 csau_3018_i406(A[3678941:3675924],A[3681959:3678942],A[3684977:3681960],tree_1[2453633:2450616],tree_1[2456651:2453634]);
csa_3018 csau_3018_i407(A[3687995:3684978],A[3691013:3687996],A[3694031:3691014],tree_1[2459669:2456652],tree_1[2462687:2459670]);
csa_3018 csau_3018_i408(A[3697049:3694032],A[3700067:3697050],A[3703085:3700068],tree_1[2465705:2462688],tree_1[2468723:2465706]);
csa_3018 csau_3018_i409(A[3706103:3703086],A[3709121:3706104],A[3712139:3709122],tree_1[2471741:2468724],tree_1[2474759:2471742]);
csa_3018 csau_3018_i410(A[3715157:3712140],A[3718175:3715158],A[3721193:3718176],tree_1[2477777:2474760],tree_1[2480795:2477778]);
csa_3018 csau_3018_i411(A[3724211:3721194],A[3727229:3724212],A[3730247:3727230],tree_1[2483813:2480796],tree_1[2486831:2483814]);
csa_3018 csau_3018_i412(A[3733265:3730248],A[3736283:3733266],A[3739301:3736284],tree_1[2489849:2486832],tree_1[2492867:2489850]);
csa_3018 csau_3018_i413(A[3742319:3739302],A[3745337:3742320],A[3748355:3745338],tree_1[2495885:2492868],tree_1[2498903:2495886]);
csa_3018 csau_3018_i414(A[3751373:3748356],A[3754391:3751374],A[3757409:3754392],tree_1[2501921:2498904],tree_1[2504939:2501922]);
csa_3018 csau_3018_i415(A[3760427:3757410],A[3763445:3760428],A[3766463:3763446],tree_1[2507957:2504940],tree_1[2510975:2507958]);
csa_3018 csau_3018_i416(A[3769481:3766464],A[3772499:3769482],A[3775517:3772500],tree_1[2513993:2510976],tree_1[2517011:2513994]);
csa_3018 csau_3018_i417(A[3778535:3775518],A[3781553:3778536],A[3784571:3781554],tree_1[2520029:2517012],tree_1[2523047:2520030]);
csa_3018 csau_3018_i418(A[3787589:3784572],A[3790607:3787590],A[3793625:3790608],tree_1[2526065:2523048],tree_1[2529083:2526066]);
csa_3018 csau_3018_i419(A[3796643:3793626],A[3799661:3796644],A[3802679:3799662],tree_1[2532101:2529084],tree_1[2535119:2532102]);
csa_3018 csau_3018_i420(A[3805697:3802680],A[3808715:3805698],A[3811733:3808716],tree_1[2538137:2535120],tree_1[2541155:2538138]);
csa_3018 csau_3018_i421(A[3814751:3811734],A[3817769:3814752],A[3820787:3817770],tree_1[2544173:2541156],tree_1[2547191:2544174]);
csa_3018 csau_3018_i422(A[3823805:3820788],A[3826823:3823806],A[3829841:3826824],tree_1[2550209:2547192],tree_1[2553227:2550210]);
csa_3018 csau_3018_i423(A[3832859:3829842],A[3835877:3832860],A[3838895:3835878],tree_1[2556245:2553228],tree_1[2559263:2556246]);
csa_3018 csau_3018_i424(A[3841913:3838896],A[3844931:3841914],A[3847949:3844932],tree_1[2562281:2559264],tree_1[2565299:2562282]);
csa_3018 csau_3018_i425(A[3850967:3847950],A[3853985:3850968],A[3857003:3853986],tree_1[2568317:2565300],tree_1[2571335:2568318]);
csa_3018 csau_3018_i426(A[3860021:3857004],A[3863039:3860022],A[3866057:3863040],tree_1[2574353:2571336],tree_1[2577371:2574354]);
csa_3018 csau_3018_i427(A[3869075:3866058],A[3872093:3869076],A[3875111:3872094],tree_1[2580389:2577372],tree_1[2583407:2580390]);
csa_3018 csau_3018_i428(A[3878129:3875112],A[3881147:3878130],A[3884165:3881148],tree_1[2586425:2583408],tree_1[2589443:2586426]);
csa_3018 csau_3018_i429(A[3887183:3884166],A[3890201:3887184],A[3893219:3890202],tree_1[2592461:2589444],tree_1[2595479:2592462]);
csa_3018 csau_3018_i430(A[3896237:3893220],A[3899255:3896238],A[3902273:3899256],tree_1[2598497:2595480],tree_1[2601515:2598498]);
csa_3018 csau_3018_i431(A[3905291:3902274],A[3908309:3905292],A[3911327:3908310],tree_1[2604533:2601516],tree_1[2607551:2604534]);
csa_3018 csau_3018_i432(A[3914345:3911328],A[3917363:3914346],A[3920381:3917364],tree_1[2610569:2607552],tree_1[2613587:2610570]);
csa_3018 csau_3018_i433(A[3923399:3920382],A[3926417:3923400],A[3929435:3926418],tree_1[2616605:2613588],tree_1[2619623:2616606]);
csa_3018 csau_3018_i434(A[3932453:3929436],A[3935471:3932454],A[3938489:3935472],tree_1[2622641:2619624],tree_1[2625659:2622642]);
csa_3018 csau_3018_i435(A[3941507:3938490],A[3944525:3941508],A[3947543:3944526],tree_1[2628677:2625660],tree_1[2631695:2628678]);
csa_3018 csau_3018_i436(A[3950561:3947544],A[3953579:3950562],A[3956597:3953580],tree_1[2634713:2631696],tree_1[2637731:2634714]);
csa_3018 csau_3018_i437(A[3959615:3956598],A[3962633:3959616],A[3965651:3962634],tree_1[2640749:2637732],tree_1[2643767:2640750]);
csa_3018 csau_3018_i438(A[3968669:3965652],A[3971687:3968670],A[3974705:3971688],tree_1[2646785:2643768],tree_1[2649803:2646786]);
csa_3018 csau_3018_i439(A[3977723:3974706],A[3980741:3977724],A[3983759:3980742],tree_1[2652821:2649804],tree_1[2655839:2652822]);
csa_3018 csau_3018_i440(A[3986777:3983760],A[3989795:3986778],A[3992813:3989796],tree_1[2658857:2655840],tree_1[2661875:2658858]);
csa_3018 csau_3018_i441(A[3995831:3992814],A[3998849:3995832],A[4001867:3998850],tree_1[2664893:2661876],tree_1[2667911:2664894]);
csa_3018 csau_3018_i442(A[4004885:4001868],A[4007903:4004886],A[4010921:4007904],tree_1[2670929:2667912],tree_1[2673947:2670930]);
csa_3018 csau_3018_i443(A[4013939:4010922],A[4016957:4013940],A[4019975:4016958],tree_1[2676965:2673948],tree_1[2679983:2676966]);
csa_3018 csau_3018_i444(A[4022993:4019976],A[4026011:4022994],A[4029029:4026012],tree_1[2683001:2679984],tree_1[2686019:2683002]);
csa_3018 csau_3018_i445(A[4032047:4029030],A[4035065:4032048],A[4038083:4035066],tree_1[2689037:2686020],tree_1[2692055:2689038]);
csa_3018 csau_3018_i446(A[4041101:4038084],A[4044119:4041102],A[4047137:4044120],tree_1[2695073:2692056],tree_1[2698091:2695074]);
csa_3018 csau_3018_i447(A[4050155:4047138],A[4053173:4050156],A[4056191:4053174],tree_1[2701109:2698092],tree_1[2704127:2701110]);
csa_3018 csau_3018_i448(A[4059209:4056192],A[4062227:4059210],A[4065245:4062228],tree_1[2707145:2704128],tree_1[2710163:2707146]);
csa_3018 csau_3018_i449(A[4068263:4065246],A[4071281:4068264],A[4074299:4071282],tree_1[2713181:2710164],tree_1[2716199:2713182]);
csa_3018 csau_3018_i450(A[4077317:4074300],A[4080335:4077318],A[4083353:4080336],tree_1[2719217:2716200],tree_1[2722235:2719218]);
csa_3018 csau_3018_i451(A[4086371:4083354],A[4089389:4086372],A[4092407:4089390],tree_1[2725253:2722236],tree_1[2728271:2725254]);
csa_3018 csau_3018_i452(A[4095425:4092408],A[4098443:4095426],A[4101461:4098444],tree_1[2731289:2728272],tree_1[2734307:2731290]);
csa_3018 csau_3018_i453(A[4104479:4101462],A[4107497:4104480],A[4110515:4107498],tree_1[2737325:2734308],tree_1[2740343:2737326]);
csa_3018 csau_3018_i454(A[4113533:4110516],A[4116551:4113534],A[4119569:4116552],tree_1[2743361:2740344],tree_1[2746379:2743362]);
csa_3018 csau_3018_i455(A[4122587:4119570],A[4125605:4122588],A[4128623:4125606],tree_1[2749397:2746380],tree_1[2752415:2749398]);
csa_3018 csau_3018_i456(A[4131641:4128624],A[4134659:4131642],A[4137677:4134660],tree_1[2755433:2752416],tree_1[2758451:2755434]);
csa_3018 csau_3018_i457(A[4140695:4137678],A[4143713:4140696],A[4146731:4143714],tree_1[2761469:2758452],tree_1[2764487:2761470]);
csa_3018 csau_3018_i458(A[4149749:4146732],A[4152767:4149750],A[4155785:4152768],tree_1[2767505:2764488],tree_1[2770523:2767506]);
csa_3018 csau_3018_i459(A[4158803:4155786],A[4161821:4158804],A[4164839:4161822],tree_1[2773541:2770524],tree_1[2776559:2773542]);
csa_3018 csau_3018_i460(A[4167857:4164840],A[4170875:4167858],A[4173893:4170876],tree_1[2779577:2776560],tree_1[2782595:2779578]);
csa_3018 csau_3018_i461(A[4176911:4173894],A[4179929:4176912],A[4182947:4179930],tree_1[2785613:2782596],tree_1[2788631:2785614]);
csa_3018 csau_3018_i462(A[4185965:4182948],A[4188983:4185966],A[4192001:4188984],tree_1[2791649:2788632],tree_1[2794667:2791650]);
csa_3018 csau_3018_i463(A[4195019:4192002],A[4198037:4195020],A[4201055:4198038],tree_1[2797685:2794668],tree_1[2800703:2797686]);
csa_3018 csau_3018_i464(A[4204073:4201056],A[4207091:4204074],A[4210109:4207092],tree_1[2803721:2800704],tree_1[2806739:2803722]);
csa_3018 csau_3018_i465(A[4213127:4210110],A[4216145:4213128],A[4219163:4216146],tree_1[2809757:2806740],tree_1[2812775:2809758]);
csa_3018 csau_3018_i466(A[4222181:4219164],A[4225199:4222182],A[4228217:4225200],tree_1[2815793:2812776],tree_1[2818811:2815794]);
csa_3018 csau_3018_i467(A[4231235:4228218],A[4234253:4231236],A[4237271:4234254],tree_1[2821829:2818812],tree_1[2824847:2821830]);
csa_3018 csau_3018_i468(A[4240289:4237272],A[4243307:4240290],A[4246325:4243308],tree_1[2827865:2824848],tree_1[2830883:2827866]);
csa_3018 csau_3018_i469(A[4249343:4246326],A[4252361:4249344],A[4255379:4252362],tree_1[2833901:2830884],tree_1[2836919:2833902]);
csa_3018 csau_3018_i470(A[4258397:4255380],A[4261415:4258398],A[4264433:4261416],tree_1[2839937:2836920],tree_1[2842955:2839938]);
csa_3018 csau_3018_i471(A[4267451:4264434],A[4270469:4267452],A[4273487:4270470],tree_1[2845973:2842956],tree_1[2848991:2845974]);
csa_3018 csau_3018_i472(A[4276505:4273488],A[4279523:4276506],A[4282541:4279524],tree_1[2852009:2848992],tree_1[2855027:2852010]);
csa_3018 csau_3018_i473(A[4285559:4282542],A[4288577:4285560],A[4291595:4288578],tree_1[2858045:2855028],tree_1[2861063:2858046]);
csa_3018 csau_3018_i474(A[4294613:4291596],A[4297631:4294614],A[4300649:4297632],tree_1[2864081:2861064],tree_1[2867099:2864082]);
csa_3018 csau_3018_i475(A[4303667:4300650],A[4306685:4303668],A[4309703:4306686],tree_1[2870117:2867100],tree_1[2873135:2870118]);
csa_3018 csau_3018_i476(A[4312721:4309704],A[4315739:4312722],A[4318757:4315740],tree_1[2876153:2873136],tree_1[2879171:2876154]);
csa_3018 csau_3018_i477(A[4321775:4318758],A[4324793:4321776],A[4327811:4324794],tree_1[2882189:2879172],tree_1[2885207:2882190]);
csa_3018 csau_3018_i478(A[4330829:4327812],A[4333847:4330830],A[4336865:4333848],tree_1[2888225:2885208],tree_1[2891243:2888226]);
csa_3018 csau_3018_i479(A[4339883:4336866],A[4342901:4339884],A[4345919:4342902],tree_1[2894261:2891244],tree_1[2897279:2894262]);
csa_3018 csau_3018_i480(A[4348937:4345920],A[4351955:4348938],A[4354973:4351956],tree_1[2900297:2897280],tree_1[2903315:2900298]);
csa_3018 csau_3018_i481(A[4357991:4354974],A[4361009:4357992],A[4364027:4361010],tree_1[2906333:2903316],tree_1[2909351:2906334]);
csa_3018 csau_3018_i482(A[4367045:4364028],A[4370063:4367046],A[4373081:4370064],tree_1[2912369:2909352],tree_1[2915387:2912370]);
csa_3018 csau_3018_i483(A[4376099:4373082],A[4379117:4376100],A[4382135:4379118],tree_1[2918405:2915388],tree_1[2921423:2918406]);
csa_3018 csau_3018_i484(A[4385153:4382136],A[4388171:4385154],A[4391189:4388172],tree_1[2924441:2921424],tree_1[2927459:2924442]);
csa_3018 csau_3018_i485(A[4394207:4391190],A[4397225:4394208],A[4400243:4397226],tree_1[2930477:2927460],tree_1[2933495:2930478]);
csa_3018 csau_3018_i486(A[4403261:4400244],A[4406279:4403262],A[4409297:4406280],tree_1[2936513:2933496],tree_1[2939531:2936514]);
csa_3018 csau_3018_i487(A[4412315:4409298],A[4415333:4412316],A[4418351:4415334],tree_1[2942549:2939532],tree_1[2945567:2942550]);
csa_3018 csau_3018_i488(A[4421369:4418352],A[4424387:4421370],A[4427405:4424388],tree_1[2948585:2945568],tree_1[2951603:2948586]);
csa_3018 csau_3018_i489(A[4430423:4427406],A[4433441:4430424],A[4436459:4433442],tree_1[2954621:2951604],tree_1[2957639:2954622]);
csa_3018 csau_3018_i490(A[4439477:4436460],A[4442495:4439478],A[4445513:4442496],tree_1[2960657:2957640],tree_1[2963675:2960658]);
csa_3018 csau_3018_i491(A[4448531:4445514],A[4451549:4448532],A[4454567:4451550],tree_1[2966693:2963676],tree_1[2969711:2966694]);
csa_3018 csau_3018_i492(A[4457585:4454568],A[4460603:4457586],A[4463621:4460604],tree_1[2972729:2969712],tree_1[2975747:2972730]);
csa_3018 csau_3018_i493(A[4466639:4463622],A[4469657:4466640],A[4472675:4469658],tree_1[2978765:2975748],tree_1[2981783:2978766]);
csa_3018 csau_3018_i494(A[4475693:4472676],A[4478711:4475694],A[4481729:4478712],tree_1[2984801:2981784],tree_1[2987819:2984802]);
csa_3018 csau_3018_i495(A[4484747:4481730],A[4487765:4484748],A[4490783:4487766],tree_1[2990837:2987820],tree_1[2993855:2990838]);
csa_3018 csau_3018_i496(A[4493801:4490784],A[4496819:4493802],A[4499837:4496820],tree_1[2996873:2993856],tree_1[2999891:2996874]);
csa_3018 csau_3018_i497(A[4502855:4499838],A[4505873:4502856],A[4508891:4505874],tree_1[3002909:2999892],tree_1[3005927:3002910]);
csa_3018 csau_3018_i498(A[4511909:4508892],A[4514927:4511910],A[4517945:4514928],tree_1[3008945:3005928],tree_1[3011963:3008946]);
csa_3018 csau_3018_i499(A[4520963:4517946],A[4523981:4520964],A[4526999:4523982],tree_1[3014981:3011964],tree_1[3017999:3014982]);
csa_3018 csau_3018_i500(A[4530017:4527000],A[4533035:4530018],A[4536053:4533036],tree_1[3021017:3018000],tree_1[3024035:3021018]);
csa_3018 csau_3018_i501(A[4539071:4536054],A[4542089:4539072],A[4545107:4542090],tree_1[3027053:3024036],tree_1[3030071:3027054]);
csa_3018 csau_3018_i502(A[4548125:4545108],A[4551143:4548126],A[4554161:4551144],tree_1[3033089:3030072],tree_1[3036107:3033090]);
// layer-2
csa_3018 csau_3018_i503(tree_1[3017:0],tree_1[6035:3018],tree_1[9053:6036],tree_2[3017:0],tree_2[6035:3018]);
csa_3018 csau_3018_i504(tree_1[12071:9054],tree_1[15089:12072],tree_1[18107:15090],tree_2[9053:6036],tree_2[12071:9054]);
csa_3018 csau_3018_i505(tree_1[21125:18108],tree_1[24143:21126],tree_1[27161:24144],tree_2[15089:12072],tree_2[18107:15090]);
csa_3018 csau_3018_i506(tree_1[30179:27162],tree_1[33197:30180],tree_1[36215:33198],tree_2[21125:18108],tree_2[24143:21126]);
csa_3018 csau_3018_i507(tree_1[39233:36216],tree_1[42251:39234],tree_1[45269:42252],tree_2[27161:24144],tree_2[30179:27162]);
csa_3018 csau_3018_i508(tree_1[48287:45270],tree_1[51305:48288],tree_1[54323:51306],tree_2[33197:30180],tree_2[36215:33198]);
csa_3018 csau_3018_i509(tree_1[57341:54324],tree_1[60359:57342],tree_1[63377:60360],tree_2[39233:36216],tree_2[42251:39234]);
csa_3018 csau_3018_i510(tree_1[66395:63378],tree_1[69413:66396],tree_1[72431:69414],tree_2[45269:42252],tree_2[48287:45270]);
csa_3018 csau_3018_i511(tree_1[75449:72432],tree_1[78467:75450],tree_1[81485:78468],tree_2[51305:48288],tree_2[54323:51306]);
csa_3018 csau_3018_i512(tree_1[84503:81486],tree_1[87521:84504],tree_1[90539:87522],tree_2[57341:54324],tree_2[60359:57342]);
csa_3018 csau_3018_i513(tree_1[93557:90540],tree_1[96575:93558],tree_1[99593:96576],tree_2[63377:60360],tree_2[66395:63378]);
csa_3018 csau_3018_i514(tree_1[102611:99594],tree_1[105629:102612],tree_1[108647:105630],tree_2[69413:66396],tree_2[72431:69414]);
csa_3018 csau_3018_i515(tree_1[111665:108648],tree_1[114683:111666],tree_1[117701:114684],tree_2[75449:72432],tree_2[78467:75450]);
csa_3018 csau_3018_i516(tree_1[120719:117702],tree_1[123737:120720],tree_1[126755:123738],tree_2[81485:78468],tree_2[84503:81486]);
csa_3018 csau_3018_i517(tree_1[129773:126756],tree_1[132791:129774],tree_1[135809:132792],tree_2[87521:84504],tree_2[90539:87522]);
csa_3018 csau_3018_i518(tree_1[138827:135810],tree_1[141845:138828],tree_1[144863:141846],tree_2[93557:90540],tree_2[96575:93558]);
csa_3018 csau_3018_i519(tree_1[147881:144864],tree_1[150899:147882],tree_1[153917:150900],tree_2[99593:96576],tree_2[102611:99594]);
csa_3018 csau_3018_i520(tree_1[156935:153918],tree_1[159953:156936],tree_1[162971:159954],tree_2[105629:102612],tree_2[108647:105630]);
csa_3018 csau_3018_i521(tree_1[165989:162972],tree_1[169007:165990],tree_1[172025:169008],tree_2[111665:108648],tree_2[114683:111666]);
csa_3018 csau_3018_i522(tree_1[175043:172026],tree_1[178061:175044],tree_1[181079:178062],tree_2[117701:114684],tree_2[120719:117702]);
csa_3018 csau_3018_i523(tree_1[184097:181080],tree_1[187115:184098],tree_1[190133:187116],tree_2[123737:120720],tree_2[126755:123738]);
csa_3018 csau_3018_i524(tree_1[193151:190134],tree_1[196169:193152],tree_1[199187:196170],tree_2[129773:126756],tree_2[132791:129774]);
csa_3018 csau_3018_i525(tree_1[202205:199188],tree_1[205223:202206],tree_1[208241:205224],tree_2[135809:132792],tree_2[138827:135810]);
csa_3018 csau_3018_i526(tree_1[211259:208242],tree_1[214277:211260],tree_1[217295:214278],tree_2[141845:138828],tree_2[144863:141846]);
csa_3018 csau_3018_i527(tree_1[220313:217296],tree_1[223331:220314],tree_1[226349:223332],tree_2[147881:144864],tree_2[150899:147882]);
csa_3018 csau_3018_i528(tree_1[229367:226350],tree_1[232385:229368],tree_1[235403:232386],tree_2[153917:150900],tree_2[156935:153918]);
csa_3018 csau_3018_i529(tree_1[238421:235404],tree_1[241439:238422],tree_1[244457:241440],tree_2[159953:156936],tree_2[162971:159954]);
csa_3018 csau_3018_i530(tree_1[247475:244458],tree_1[250493:247476],tree_1[253511:250494],tree_2[165989:162972],tree_2[169007:165990]);
csa_3018 csau_3018_i531(tree_1[256529:253512],tree_1[259547:256530],tree_1[262565:259548],tree_2[172025:169008],tree_2[175043:172026]);
csa_3018 csau_3018_i532(tree_1[265583:262566],tree_1[268601:265584],tree_1[271619:268602],tree_2[178061:175044],tree_2[181079:178062]);
csa_3018 csau_3018_i533(tree_1[274637:271620],tree_1[277655:274638],tree_1[280673:277656],tree_2[184097:181080],tree_2[187115:184098]);
csa_3018 csau_3018_i534(tree_1[283691:280674],tree_1[286709:283692],tree_1[289727:286710],tree_2[190133:187116],tree_2[193151:190134]);
csa_3018 csau_3018_i535(tree_1[292745:289728],tree_1[295763:292746],tree_1[298781:295764],tree_2[196169:193152],tree_2[199187:196170]);
csa_3018 csau_3018_i536(tree_1[301799:298782],tree_1[304817:301800],tree_1[307835:304818],tree_2[202205:199188],tree_2[205223:202206]);
csa_3018 csau_3018_i537(tree_1[310853:307836],tree_1[313871:310854],tree_1[316889:313872],tree_2[208241:205224],tree_2[211259:208242]);
csa_3018 csau_3018_i538(tree_1[319907:316890],tree_1[322925:319908],tree_1[325943:322926],tree_2[214277:211260],tree_2[217295:214278]);
csa_3018 csau_3018_i539(tree_1[328961:325944],tree_1[331979:328962],tree_1[334997:331980],tree_2[220313:217296],tree_2[223331:220314]);
csa_3018 csau_3018_i540(tree_1[338015:334998],tree_1[341033:338016],tree_1[344051:341034],tree_2[226349:223332],tree_2[229367:226350]);
csa_3018 csau_3018_i541(tree_1[347069:344052],tree_1[350087:347070],tree_1[353105:350088],tree_2[232385:229368],tree_2[235403:232386]);
csa_3018 csau_3018_i542(tree_1[356123:353106],tree_1[359141:356124],tree_1[362159:359142],tree_2[238421:235404],tree_2[241439:238422]);
csa_3018 csau_3018_i543(tree_1[365177:362160],tree_1[368195:365178],tree_1[371213:368196],tree_2[244457:241440],tree_2[247475:244458]);
csa_3018 csau_3018_i544(tree_1[374231:371214],tree_1[377249:374232],tree_1[380267:377250],tree_2[250493:247476],tree_2[253511:250494]);
csa_3018 csau_3018_i545(tree_1[383285:380268],tree_1[386303:383286],tree_1[389321:386304],tree_2[256529:253512],tree_2[259547:256530]);
csa_3018 csau_3018_i546(tree_1[392339:389322],tree_1[395357:392340],tree_1[398375:395358],tree_2[262565:259548],tree_2[265583:262566]);
csa_3018 csau_3018_i547(tree_1[401393:398376],tree_1[404411:401394],tree_1[407429:404412],tree_2[268601:265584],tree_2[271619:268602]);
csa_3018 csau_3018_i548(tree_1[410447:407430],tree_1[413465:410448],tree_1[416483:413466],tree_2[274637:271620],tree_2[277655:274638]);
csa_3018 csau_3018_i549(tree_1[419501:416484],tree_1[422519:419502],tree_1[425537:422520],tree_2[280673:277656],tree_2[283691:280674]);
csa_3018 csau_3018_i550(tree_1[428555:425538],tree_1[431573:428556],tree_1[434591:431574],tree_2[286709:283692],tree_2[289727:286710]);
csa_3018 csau_3018_i551(tree_1[437609:434592],tree_1[440627:437610],tree_1[443645:440628],tree_2[292745:289728],tree_2[295763:292746]);
csa_3018 csau_3018_i552(tree_1[446663:443646],tree_1[449681:446664],tree_1[452699:449682],tree_2[298781:295764],tree_2[301799:298782]);
csa_3018 csau_3018_i553(tree_1[455717:452700],tree_1[458735:455718],tree_1[461753:458736],tree_2[304817:301800],tree_2[307835:304818]);
csa_3018 csau_3018_i554(tree_1[464771:461754],tree_1[467789:464772],tree_1[470807:467790],tree_2[310853:307836],tree_2[313871:310854]);
csa_3018 csau_3018_i555(tree_1[473825:470808],tree_1[476843:473826],tree_1[479861:476844],tree_2[316889:313872],tree_2[319907:316890]);
csa_3018 csau_3018_i556(tree_1[482879:479862],tree_1[485897:482880],tree_1[488915:485898],tree_2[322925:319908],tree_2[325943:322926]);
csa_3018 csau_3018_i557(tree_1[491933:488916],tree_1[494951:491934],tree_1[497969:494952],tree_2[328961:325944],tree_2[331979:328962]);
csa_3018 csau_3018_i558(tree_1[500987:497970],tree_1[504005:500988],tree_1[507023:504006],tree_2[334997:331980],tree_2[338015:334998]);
csa_3018 csau_3018_i559(tree_1[510041:507024],tree_1[513059:510042],tree_1[516077:513060],tree_2[341033:338016],tree_2[344051:341034]);
csa_3018 csau_3018_i560(tree_1[519095:516078],tree_1[522113:519096],tree_1[525131:522114],tree_2[347069:344052],tree_2[350087:347070]);
csa_3018 csau_3018_i561(tree_1[528149:525132],tree_1[531167:528150],tree_1[534185:531168],tree_2[353105:350088],tree_2[356123:353106]);
csa_3018 csau_3018_i562(tree_1[537203:534186],tree_1[540221:537204],tree_1[543239:540222],tree_2[359141:356124],tree_2[362159:359142]);
csa_3018 csau_3018_i563(tree_1[546257:543240],tree_1[549275:546258],tree_1[552293:549276],tree_2[365177:362160],tree_2[368195:365178]);
csa_3018 csau_3018_i564(tree_1[555311:552294],tree_1[558329:555312],tree_1[561347:558330],tree_2[371213:368196],tree_2[374231:371214]);
csa_3018 csau_3018_i565(tree_1[564365:561348],tree_1[567383:564366],tree_1[570401:567384],tree_2[377249:374232],tree_2[380267:377250]);
csa_3018 csau_3018_i566(tree_1[573419:570402],tree_1[576437:573420],tree_1[579455:576438],tree_2[383285:380268],tree_2[386303:383286]);
csa_3018 csau_3018_i567(tree_1[582473:579456],tree_1[585491:582474],tree_1[588509:585492],tree_2[389321:386304],tree_2[392339:389322]);
csa_3018 csau_3018_i568(tree_1[591527:588510],tree_1[594545:591528],tree_1[597563:594546],tree_2[395357:392340],tree_2[398375:395358]);
csa_3018 csau_3018_i569(tree_1[600581:597564],tree_1[603599:600582],tree_1[606617:603600],tree_2[401393:398376],tree_2[404411:401394]);
csa_3018 csau_3018_i570(tree_1[609635:606618],tree_1[612653:609636],tree_1[615671:612654],tree_2[407429:404412],tree_2[410447:407430]);
csa_3018 csau_3018_i571(tree_1[618689:615672],tree_1[621707:618690],tree_1[624725:621708],tree_2[413465:410448],tree_2[416483:413466]);
csa_3018 csau_3018_i572(tree_1[627743:624726],tree_1[630761:627744],tree_1[633779:630762],tree_2[419501:416484],tree_2[422519:419502]);
csa_3018 csau_3018_i573(tree_1[636797:633780],tree_1[639815:636798],tree_1[642833:639816],tree_2[425537:422520],tree_2[428555:425538]);
csa_3018 csau_3018_i574(tree_1[645851:642834],tree_1[648869:645852],tree_1[651887:648870],tree_2[431573:428556],tree_2[434591:431574]);
csa_3018 csau_3018_i575(tree_1[654905:651888],tree_1[657923:654906],tree_1[660941:657924],tree_2[437609:434592],tree_2[440627:437610]);
csa_3018 csau_3018_i576(tree_1[663959:660942],tree_1[666977:663960],tree_1[669995:666978],tree_2[443645:440628],tree_2[446663:443646]);
csa_3018 csau_3018_i577(tree_1[673013:669996],tree_1[676031:673014],tree_1[679049:676032],tree_2[449681:446664],tree_2[452699:449682]);
csa_3018 csau_3018_i578(tree_1[682067:679050],tree_1[685085:682068],tree_1[688103:685086],tree_2[455717:452700],tree_2[458735:455718]);
csa_3018 csau_3018_i579(tree_1[691121:688104],tree_1[694139:691122],tree_1[697157:694140],tree_2[461753:458736],tree_2[464771:461754]);
csa_3018 csau_3018_i580(tree_1[700175:697158],tree_1[703193:700176],tree_1[706211:703194],tree_2[467789:464772],tree_2[470807:467790]);
csa_3018 csau_3018_i581(tree_1[709229:706212],tree_1[712247:709230],tree_1[715265:712248],tree_2[473825:470808],tree_2[476843:473826]);
csa_3018 csau_3018_i582(tree_1[718283:715266],tree_1[721301:718284],tree_1[724319:721302],tree_2[479861:476844],tree_2[482879:479862]);
csa_3018 csau_3018_i583(tree_1[727337:724320],tree_1[730355:727338],tree_1[733373:730356],tree_2[485897:482880],tree_2[488915:485898]);
csa_3018 csau_3018_i584(tree_1[736391:733374],tree_1[739409:736392],tree_1[742427:739410],tree_2[491933:488916],tree_2[494951:491934]);
csa_3018 csau_3018_i585(tree_1[745445:742428],tree_1[748463:745446],tree_1[751481:748464],tree_2[497969:494952],tree_2[500987:497970]);
csa_3018 csau_3018_i586(tree_1[754499:751482],tree_1[757517:754500],tree_1[760535:757518],tree_2[504005:500988],tree_2[507023:504006]);
csa_3018 csau_3018_i587(tree_1[763553:760536],tree_1[766571:763554],tree_1[769589:766572],tree_2[510041:507024],tree_2[513059:510042]);
csa_3018 csau_3018_i588(tree_1[772607:769590],tree_1[775625:772608],tree_1[778643:775626],tree_2[516077:513060],tree_2[519095:516078]);
csa_3018 csau_3018_i589(tree_1[781661:778644],tree_1[784679:781662],tree_1[787697:784680],tree_2[522113:519096],tree_2[525131:522114]);
csa_3018 csau_3018_i590(tree_1[790715:787698],tree_1[793733:790716],tree_1[796751:793734],tree_2[528149:525132],tree_2[531167:528150]);
csa_3018 csau_3018_i591(tree_1[799769:796752],tree_1[802787:799770],tree_1[805805:802788],tree_2[534185:531168],tree_2[537203:534186]);
csa_3018 csau_3018_i592(tree_1[808823:805806],tree_1[811841:808824],tree_1[814859:811842],tree_2[540221:537204],tree_2[543239:540222]);
csa_3018 csau_3018_i593(tree_1[817877:814860],tree_1[820895:817878],tree_1[823913:820896],tree_2[546257:543240],tree_2[549275:546258]);
csa_3018 csau_3018_i594(tree_1[826931:823914],tree_1[829949:826932],tree_1[832967:829950],tree_2[552293:549276],tree_2[555311:552294]);
csa_3018 csau_3018_i595(tree_1[835985:832968],tree_1[839003:835986],tree_1[842021:839004],tree_2[558329:555312],tree_2[561347:558330]);
csa_3018 csau_3018_i596(tree_1[845039:842022],tree_1[848057:845040],tree_1[851075:848058],tree_2[564365:561348],tree_2[567383:564366]);
csa_3018 csau_3018_i597(tree_1[854093:851076],tree_1[857111:854094],tree_1[860129:857112],tree_2[570401:567384],tree_2[573419:570402]);
csa_3018 csau_3018_i598(tree_1[863147:860130],tree_1[866165:863148],tree_1[869183:866166],tree_2[576437:573420],tree_2[579455:576438]);
csa_3018 csau_3018_i599(tree_1[872201:869184],tree_1[875219:872202],tree_1[878237:875220],tree_2[582473:579456],tree_2[585491:582474]);
csa_3018 csau_3018_i600(tree_1[881255:878238],tree_1[884273:881256],tree_1[887291:884274],tree_2[588509:585492],tree_2[591527:588510]);
csa_3018 csau_3018_i601(tree_1[890309:887292],tree_1[893327:890310],tree_1[896345:893328],tree_2[594545:591528],tree_2[597563:594546]);
csa_3018 csau_3018_i602(tree_1[899363:896346],tree_1[902381:899364],tree_1[905399:902382],tree_2[600581:597564],tree_2[603599:600582]);
csa_3018 csau_3018_i603(tree_1[908417:905400],tree_1[911435:908418],tree_1[914453:911436],tree_2[606617:603600],tree_2[609635:606618]);
csa_3018 csau_3018_i604(tree_1[917471:914454],tree_1[920489:917472],tree_1[923507:920490],tree_2[612653:609636],tree_2[615671:612654]);
csa_3018 csau_3018_i605(tree_1[926525:923508],tree_1[929543:926526],tree_1[932561:929544],tree_2[618689:615672],tree_2[621707:618690]);
csa_3018 csau_3018_i606(tree_1[935579:932562],tree_1[938597:935580],tree_1[941615:938598],tree_2[624725:621708],tree_2[627743:624726]);
csa_3018 csau_3018_i607(tree_1[944633:941616],tree_1[947651:944634],tree_1[950669:947652],tree_2[630761:627744],tree_2[633779:630762]);
csa_3018 csau_3018_i608(tree_1[953687:950670],tree_1[956705:953688],tree_1[959723:956706],tree_2[636797:633780],tree_2[639815:636798]);
csa_3018 csau_3018_i609(tree_1[962741:959724],tree_1[965759:962742],tree_1[968777:965760],tree_2[642833:639816],tree_2[645851:642834]);
csa_3018 csau_3018_i610(tree_1[971795:968778],tree_1[974813:971796],tree_1[977831:974814],tree_2[648869:645852],tree_2[651887:648870]);
csa_3018 csau_3018_i611(tree_1[980849:977832],tree_1[983867:980850],tree_1[986885:983868],tree_2[654905:651888],tree_2[657923:654906]);
csa_3018 csau_3018_i612(tree_1[989903:986886],tree_1[992921:989904],tree_1[995939:992922],tree_2[660941:657924],tree_2[663959:660942]);
csa_3018 csau_3018_i613(tree_1[998957:995940],tree_1[1001975:998958],tree_1[1004993:1001976],tree_2[666977:663960],tree_2[669995:666978]);
csa_3018 csau_3018_i614(tree_1[1008011:1004994],tree_1[1011029:1008012],tree_1[1014047:1011030],tree_2[673013:669996],tree_2[676031:673014]);
csa_3018 csau_3018_i615(tree_1[1017065:1014048],tree_1[1020083:1017066],tree_1[1023101:1020084],tree_2[679049:676032],tree_2[682067:679050]);
csa_3018 csau_3018_i616(tree_1[1026119:1023102],tree_1[1029137:1026120],tree_1[1032155:1029138],tree_2[685085:682068],tree_2[688103:685086]);
csa_3018 csau_3018_i617(tree_1[1035173:1032156],tree_1[1038191:1035174],tree_1[1041209:1038192],tree_2[691121:688104],tree_2[694139:691122]);
csa_3018 csau_3018_i618(tree_1[1044227:1041210],tree_1[1047245:1044228],tree_1[1050263:1047246],tree_2[697157:694140],tree_2[700175:697158]);
csa_3018 csau_3018_i619(tree_1[1053281:1050264],tree_1[1056299:1053282],tree_1[1059317:1056300],tree_2[703193:700176],tree_2[706211:703194]);
csa_3018 csau_3018_i620(tree_1[1062335:1059318],tree_1[1065353:1062336],tree_1[1068371:1065354],tree_2[709229:706212],tree_2[712247:709230]);
csa_3018 csau_3018_i621(tree_1[1071389:1068372],tree_1[1074407:1071390],tree_1[1077425:1074408],tree_2[715265:712248],tree_2[718283:715266]);
csa_3018 csau_3018_i622(tree_1[1080443:1077426],tree_1[1083461:1080444],tree_1[1086479:1083462],tree_2[721301:718284],tree_2[724319:721302]);
csa_3018 csau_3018_i623(tree_1[1089497:1086480],tree_1[1092515:1089498],tree_1[1095533:1092516],tree_2[727337:724320],tree_2[730355:727338]);
csa_3018 csau_3018_i624(tree_1[1098551:1095534],tree_1[1101569:1098552],tree_1[1104587:1101570],tree_2[733373:730356],tree_2[736391:733374]);
csa_3018 csau_3018_i625(tree_1[1107605:1104588],tree_1[1110623:1107606],tree_1[1113641:1110624],tree_2[739409:736392],tree_2[742427:739410]);
csa_3018 csau_3018_i626(tree_1[1116659:1113642],tree_1[1119677:1116660],tree_1[1122695:1119678],tree_2[745445:742428],tree_2[748463:745446]);
csa_3018 csau_3018_i627(tree_1[1125713:1122696],tree_1[1128731:1125714],tree_1[1131749:1128732],tree_2[751481:748464],tree_2[754499:751482]);
csa_3018 csau_3018_i628(tree_1[1134767:1131750],tree_1[1137785:1134768],tree_1[1140803:1137786],tree_2[757517:754500],tree_2[760535:757518]);
csa_3018 csau_3018_i629(tree_1[1143821:1140804],tree_1[1146839:1143822],tree_1[1149857:1146840],tree_2[763553:760536],tree_2[766571:763554]);
csa_3018 csau_3018_i630(tree_1[1152875:1149858],tree_1[1155893:1152876],tree_1[1158911:1155894],tree_2[769589:766572],tree_2[772607:769590]);
csa_3018 csau_3018_i631(tree_1[1161929:1158912],tree_1[1164947:1161930],tree_1[1167965:1164948],tree_2[775625:772608],tree_2[778643:775626]);
csa_3018 csau_3018_i632(tree_1[1170983:1167966],tree_1[1174001:1170984],tree_1[1177019:1174002],tree_2[781661:778644],tree_2[784679:781662]);
csa_3018 csau_3018_i633(tree_1[1180037:1177020],tree_1[1183055:1180038],tree_1[1186073:1183056],tree_2[787697:784680],tree_2[790715:787698]);
csa_3018 csau_3018_i634(tree_1[1189091:1186074],tree_1[1192109:1189092],tree_1[1195127:1192110],tree_2[793733:790716],tree_2[796751:793734]);
csa_3018 csau_3018_i635(tree_1[1198145:1195128],tree_1[1201163:1198146],tree_1[1204181:1201164],tree_2[799769:796752],tree_2[802787:799770]);
csa_3018 csau_3018_i636(tree_1[1207199:1204182],tree_1[1210217:1207200],tree_1[1213235:1210218],tree_2[805805:802788],tree_2[808823:805806]);
csa_3018 csau_3018_i637(tree_1[1216253:1213236],tree_1[1219271:1216254],tree_1[1222289:1219272],tree_2[811841:808824],tree_2[814859:811842]);
csa_3018 csau_3018_i638(tree_1[1225307:1222290],tree_1[1228325:1225308],tree_1[1231343:1228326],tree_2[817877:814860],tree_2[820895:817878]);
csa_3018 csau_3018_i639(tree_1[1234361:1231344],tree_1[1237379:1234362],tree_1[1240397:1237380],tree_2[823913:820896],tree_2[826931:823914]);
csa_3018 csau_3018_i640(tree_1[1243415:1240398],tree_1[1246433:1243416],tree_1[1249451:1246434],tree_2[829949:826932],tree_2[832967:829950]);
csa_3018 csau_3018_i641(tree_1[1252469:1249452],tree_1[1255487:1252470],tree_1[1258505:1255488],tree_2[835985:832968],tree_2[839003:835986]);
csa_3018 csau_3018_i642(tree_1[1261523:1258506],tree_1[1264541:1261524],tree_1[1267559:1264542],tree_2[842021:839004],tree_2[845039:842022]);
csa_3018 csau_3018_i643(tree_1[1270577:1267560],tree_1[1273595:1270578],tree_1[1276613:1273596],tree_2[848057:845040],tree_2[851075:848058]);
csa_3018 csau_3018_i644(tree_1[1279631:1276614],tree_1[1282649:1279632],tree_1[1285667:1282650],tree_2[854093:851076],tree_2[857111:854094]);
csa_3018 csau_3018_i645(tree_1[1288685:1285668],tree_1[1291703:1288686],tree_1[1294721:1291704],tree_2[860129:857112],tree_2[863147:860130]);
csa_3018 csau_3018_i646(tree_1[1297739:1294722],tree_1[1300757:1297740],tree_1[1303775:1300758],tree_2[866165:863148],tree_2[869183:866166]);
csa_3018 csau_3018_i647(tree_1[1306793:1303776],tree_1[1309811:1306794],tree_1[1312829:1309812],tree_2[872201:869184],tree_2[875219:872202]);
csa_3018 csau_3018_i648(tree_1[1315847:1312830],tree_1[1318865:1315848],tree_1[1321883:1318866],tree_2[878237:875220],tree_2[881255:878238]);
csa_3018 csau_3018_i649(tree_1[1324901:1321884],tree_1[1327919:1324902],tree_1[1330937:1327920],tree_2[884273:881256],tree_2[887291:884274]);
csa_3018 csau_3018_i650(tree_1[1333955:1330938],tree_1[1336973:1333956],tree_1[1339991:1336974],tree_2[890309:887292],tree_2[893327:890310]);
csa_3018 csau_3018_i651(tree_1[1343009:1339992],tree_1[1346027:1343010],tree_1[1349045:1346028],tree_2[896345:893328],tree_2[899363:896346]);
csa_3018 csau_3018_i652(tree_1[1352063:1349046],tree_1[1355081:1352064],tree_1[1358099:1355082],tree_2[902381:899364],tree_2[905399:902382]);
csa_3018 csau_3018_i653(tree_1[1361117:1358100],tree_1[1364135:1361118],tree_1[1367153:1364136],tree_2[908417:905400],tree_2[911435:908418]);
csa_3018 csau_3018_i654(tree_1[1370171:1367154],tree_1[1373189:1370172],tree_1[1376207:1373190],tree_2[914453:911436],tree_2[917471:914454]);
csa_3018 csau_3018_i655(tree_1[1379225:1376208],tree_1[1382243:1379226],tree_1[1385261:1382244],tree_2[920489:917472],tree_2[923507:920490]);
csa_3018 csau_3018_i656(tree_1[1388279:1385262],tree_1[1391297:1388280],tree_1[1394315:1391298],tree_2[926525:923508],tree_2[929543:926526]);
csa_3018 csau_3018_i657(tree_1[1397333:1394316],tree_1[1400351:1397334],tree_1[1403369:1400352],tree_2[932561:929544],tree_2[935579:932562]);
csa_3018 csau_3018_i658(tree_1[1406387:1403370],tree_1[1409405:1406388],tree_1[1412423:1409406],tree_2[938597:935580],tree_2[941615:938598]);
csa_3018 csau_3018_i659(tree_1[1415441:1412424],tree_1[1418459:1415442],tree_1[1421477:1418460],tree_2[944633:941616],tree_2[947651:944634]);
csa_3018 csau_3018_i660(tree_1[1424495:1421478],tree_1[1427513:1424496],tree_1[1430531:1427514],tree_2[950669:947652],tree_2[953687:950670]);
csa_3018 csau_3018_i661(tree_1[1433549:1430532],tree_1[1436567:1433550],tree_1[1439585:1436568],tree_2[956705:953688],tree_2[959723:956706]);
csa_3018 csau_3018_i662(tree_1[1442603:1439586],tree_1[1445621:1442604],tree_1[1448639:1445622],tree_2[962741:959724],tree_2[965759:962742]);
csa_3018 csau_3018_i663(tree_1[1451657:1448640],tree_1[1454675:1451658],tree_1[1457693:1454676],tree_2[968777:965760],tree_2[971795:968778]);
csa_3018 csau_3018_i664(tree_1[1460711:1457694],tree_1[1463729:1460712],tree_1[1466747:1463730],tree_2[974813:971796],tree_2[977831:974814]);
csa_3018 csau_3018_i665(tree_1[1469765:1466748],tree_1[1472783:1469766],tree_1[1475801:1472784],tree_2[980849:977832],tree_2[983867:980850]);
csa_3018 csau_3018_i666(tree_1[1478819:1475802],tree_1[1481837:1478820],tree_1[1484855:1481838],tree_2[986885:983868],tree_2[989903:986886]);
csa_3018 csau_3018_i667(tree_1[1487873:1484856],tree_1[1490891:1487874],tree_1[1493909:1490892],tree_2[992921:989904],tree_2[995939:992922]);
csa_3018 csau_3018_i668(tree_1[1496927:1493910],tree_1[1499945:1496928],tree_1[1502963:1499946],tree_2[998957:995940],tree_2[1001975:998958]);
csa_3018 csau_3018_i669(tree_1[1505981:1502964],tree_1[1508999:1505982],tree_1[1512017:1509000],tree_2[1004993:1001976],tree_2[1008011:1004994]);
csa_3018 csau_3018_i670(tree_1[1515035:1512018],tree_1[1518053:1515036],tree_1[1521071:1518054],tree_2[1011029:1008012],tree_2[1014047:1011030]);
csa_3018 csau_3018_i671(tree_1[1524089:1521072],tree_1[1527107:1524090],tree_1[1530125:1527108],tree_2[1017065:1014048],tree_2[1020083:1017066]);
csa_3018 csau_3018_i672(tree_1[1533143:1530126],tree_1[1536161:1533144],tree_1[1539179:1536162],tree_2[1023101:1020084],tree_2[1026119:1023102]);
csa_3018 csau_3018_i673(tree_1[1542197:1539180],tree_1[1545215:1542198],tree_1[1548233:1545216],tree_2[1029137:1026120],tree_2[1032155:1029138]);
csa_3018 csau_3018_i674(tree_1[1551251:1548234],tree_1[1554269:1551252],tree_1[1557287:1554270],tree_2[1035173:1032156],tree_2[1038191:1035174]);
csa_3018 csau_3018_i675(tree_1[1560305:1557288],tree_1[1563323:1560306],tree_1[1566341:1563324],tree_2[1041209:1038192],tree_2[1044227:1041210]);
csa_3018 csau_3018_i676(tree_1[1569359:1566342],tree_1[1572377:1569360],tree_1[1575395:1572378],tree_2[1047245:1044228],tree_2[1050263:1047246]);
csa_3018 csau_3018_i677(tree_1[1578413:1575396],tree_1[1581431:1578414],tree_1[1584449:1581432],tree_2[1053281:1050264],tree_2[1056299:1053282]);
csa_3018 csau_3018_i678(tree_1[1587467:1584450],tree_1[1590485:1587468],tree_1[1593503:1590486],tree_2[1059317:1056300],tree_2[1062335:1059318]);
csa_3018 csau_3018_i679(tree_1[1596521:1593504],tree_1[1599539:1596522],tree_1[1602557:1599540],tree_2[1065353:1062336],tree_2[1068371:1065354]);
csa_3018 csau_3018_i680(tree_1[1605575:1602558],tree_1[1608593:1605576],tree_1[1611611:1608594],tree_2[1071389:1068372],tree_2[1074407:1071390]);
csa_3018 csau_3018_i681(tree_1[1614629:1611612],tree_1[1617647:1614630],tree_1[1620665:1617648],tree_2[1077425:1074408],tree_2[1080443:1077426]);
csa_3018 csau_3018_i682(tree_1[1623683:1620666],tree_1[1626701:1623684],tree_1[1629719:1626702],tree_2[1083461:1080444],tree_2[1086479:1083462]);
csa_3018 csau_3018_i683(tree_1[1632737:1629720],tree_1[1635755:1632738],tree_1[1638773:1635756],tree_2[1089497:1086480],tree_2[1092515:1089498]);
csa_3018 csau_3018_i684(tree_1[1641791:1638774],tree_1[1644809:1641792],tree_1[1647827:1644810],tree_2[1095533:1092516],tree_2[1098551:1095534]);
csa_3018 csau_3018_i685(tree_1[1650845:1647828],tree_1[1653863:1650846],tree_1[1656881:1653864],tree_2[1101569:1098552],tree_2[1104587:1101570]);
csa_3018 csau_3018_i686(tree_1[1659899:1656882],tree_1[1662917:1659900],tree_1[1665935:1662918],tree_2[1107605:1104588],tree_2[1110623:1107606]);
csa_3018 csau_3018_i687(tree_1[1668953:1665936],tree_1[1671971:1668954],tree_1[1674989:1671972],tree_2[1113641:1110624],tree_2[1116659:1113642]);
csa_3018 csau_3018_i688(tree_1[1678007:1674990],tree_1[1681025:1678008],tree_1[1684043:1681026],tree_2[1119677:1116660],tree_2[1122695:1119678]);
csa_3018 csau_3018_i689(tree_1[1687061:1684044],tree_1[1690079:1687062],tree_1[1693097:1690080],tree_2[1125713:1122696],tree_2[1128731:1125714]);
csa_3018 csau_3018_i690(tree_1[1696115:1693098],tree_1[1699133:1696116],tree_1[1702151:1699134],tree_2[1131749:1128732],tree_2[1134767:1131750]);
csa_3018 csau_3018_i691(tree_1[1705169:1702152],tree_1[1708187:1705170],tree_1[1711205:1708188],tree_2[1137785:1134768],tree_2[1140803:1137786]);
csa_3018 csau_3018_i692(tree_1[1714223:1711206],tree_1[1717241:1714224],tree_1[1720259:1717242],tree_2[1143821:1140804],tree_2[1146839:1143822]);
csa_3018 csau_3018_i693(tree_1[1723277:1720260],tree_1[1726295:1723278],tree_1[1729313:1726296],tree_2[1149857:1146840],tree_2[1152875:1149858]);
csa_3018 csau_3018_i694(tree_1[1732331:1729314],tree_1[1735349:1732332],tree_1[1738367:1735350],tree_2[1155893:1152876],tree_2[1158911:1155894]);
csa_3018 csau_3018_i695(tree_1[1741385:1738368],tree_1[1744403:1741386],tree_1[1747421:1744404],tree_2[1161929:1158912],tree_2[1164947:1161930]);
csa_3018 csau_3018_i696(tree_1[1750439:1747422],tree_1[1753457:1750440],tree_1[1756475:1753458],tree_2[1167965:1164948],tree_2[1170983:1167966]);
csa_3018 csau_3018_i697(tree_1[1759493:1756476],tree_1[1762511:1759494],tree_1[1765529:1762512],tree_2[1174001:1170984],tree_2[1177019:1174002]);
csa_3018 csau_3018_i698(tree_1[1768547:1765530],tree_1[1771565:1768548],tree_1[1774583:1771566],tree_2[1180037:1177020],tree_2[1183055:1180038]);
csa_3018 csau_3018_i699(tree_1[1777601:1774584],tree_1[1780619:1777602],tree_1[1783637:1780620],tree_2[1186073:1183056],tree_2[1189091:1186074]);
csa_3018 csau_3018_i700(tree_1[1786655:1783638],tree_1[1789673:1786656],tree_1[1792691:1789674],tree_2[1192109:1189092],tree_2[1195127:1192110]);
csa_3018 csau_3018_i701(tree_1[1795709:1792692],tree_1[1798727:1795710],tree_1[1801745:1798728],tree_2[1198145:1195128],tree_2[1201163:1198146]);
csa_3018 csau_3018_i702(tree_1[1804763:1801746],tree_1[1807781:1804764],tree_1[1810799:1807782],tree_2[1204181:1201164],tree_2[1207199:1204182]);
csa_3018 csau_3018_i703(tree_1[1813817:1810800],tree_1[1816835:1813818],tree_1[1819853:1816836],tree_2[1210217:1207200],tree_2[1213235:1210218]);
csa_3018 csau_3018_i704(tree_1[1822871:1819854],tree_1[1825889:1822872],tree_1[1828907:1825890],tree_2[1216253:1213236],tree_2[1219271:1216254]);
csa_3018 csau_3018_i705(tree_1[1831925:1828908],tree_1[1834943:1831926],tree_1[1837961:1834944],tree_2[1222289:1219272],tree_2[1225307:1222290]);
csa_3018 csau_3018_i706(tree_1[1840979:1837962],tree_1[1843997:1840980],tree_1[1847015:1843998],tree_2[1228325:1225308],tree_2[1231343:1228326]);
csa_3018 csau_3018_i707(tree_1[1850033:1847016],tree_1[1853051:1850034],tree_1[1856069:1853052],tree_2[1234361:1231344],tree_2[1237379:1234362]);
csa_3018 csau_3018_i708(tree_1[1859087:1856070],tree_1[1862105:1859088],tree_1[1865123:1862106],tree_2[1240397:1237380],tree_2[1243415:1240398]);
csa_3018 csau_3018_i709(tree_1[1868141:1865124],tree_1[1871159:1868142],tree_1[1874177:1871160],tree_2[1246433:1243416],tree_2[1249451:1246434]);
csa_3018 csau_3018_i710(tree_1[1877195:1874178],tree_1[1880213:1877196],tree_1[1883231:1880214],tree_2[1252469:1249452],tree_2[1255487:1252470]);
csa_3018 csau_3018_i711(tree_1[1886249:1883232],tree_1[1889267:1886250],tree_1[1892285:1889268],tree_2[1258505:1255488],tree_2[1261523:1258506]);
csa_3018 csau_3018_i712(tree_1[1895303:1892286],tree_1[1898321:1895304],tree_1[1901339:1898322],tree_2[1264541:1261524],tree_2[1267559:1264542]);
csa_3018 csau_3018_i713(tree_1[1904357:1901340],tree_1[1907375:1904358],tree_1[1910393:1907376],tree_2[1270577:1267560],tree_2[1273595:1270578]);
csa_3018 csau_3018_i714(tree_1[1913411:1910394],tree_1[1916429:1913412],tree_1[1919447:1916430],tree_2[1276613:1273596],tree_2[1279631:1276614]);
csa_3018 csau_3018_i715(tree_1[1922465:1919448],tree_1[1925483:1922466],tree_1[1928501:1925484],tree_2[1282649:1279632],tree_2[1285667:1282650]);
csa_3018 csau_3018_i716(tree_1[1931519:1928502],tree_1[1934537:1931520],tree_1[1937555:1934538],tree_2[1288685:1285668],tree_2[1291703:1288686]);
csa_3018 csau_3018_i717(tree_1[1940573:1937556],tree_1[1943591:1940574],tree_1[1946609:1943592],tree_2[1294721:1291704],tree_2[1297739:1294722]);
csa_3018 csau_3018_i718(tree_1[1949627:1946610],tree_1[1952645:1949628],tree_1[1955663:1952646],tree_2[1300757:1297740],tree_2[1303775:1300758]);
csa_3018 csau_3018_i719(tree_1[1958681:1955664],tree_1[1961699:1958682],tree_1[1964717:1961700],tree_2[1306793:1303776],tree_2[1309811:1306794]);
csa_3018 csau_3018_i720(tree_1[1967735:1964718],tree_1[1970753:1967736],tree_1[1973771:1970754],tree_2[1312829:1309812],tree_2[1315847:1312830]);
csa_3018 csau_3018_i721(tree_1[1976789:1973772],tree_1[1979807:1976790],tree_1[1982825:1979808],tree_2[1318865:1315848],tree_2[1321883:1318866]);
csa_3018 csau_3018_i722(tree_1[1985843:1982826],tree_1[1988861:1985844],tree_1[1991879:1988862],tree_2[1324901:1321884],tree_2[1327919:1324902]);
csa_3018 csau_3018_i723(tree_1[1994897:1991880],tree_1[1997915:1994898],tree_1[2000933:1997916],tree_2[1330937:1327920],tree_2[1333955:1330938]);
csa_3018 csau_3018_i724(tree_1[2003951:2000934],tree_1[2006969:2003952],tree_1[2009987:2006970],tree_2[1336973:1333956],tree_2[1339991:1336974]);
csa_3018 csau_3018_i725(tree_1[2013005:2009988],tree_1[2016023:2013006],tree_1[2019041:2016024],tree_2[1343009:1339992],tree_2[1346027:1343010]);
csa_3018 csau_3018_i726(tree_1[2022059:2019042],tree_1[2025077:2022060],tree_1[2028095:2025078],tree_2[1349045:1346028],tree_2[1352063:1349046]);
csa_3018 csau_3018_i727(tree_1[2031113:2028096],tree_1[2034131:2031114],tree_1[2037149:2034132],tree_2[1355081:1352064],tree_2[1358099:1355082]);
csa_3018 csau_3018_i728(tree_1[2040167:2037150],tree_1[2043185:2040168],tree_1[2046203:2043186],tree_2[1361117:1358100],tree_2[1364135:1361118]);
csa_3018 csau_3018_i729(tree_1[2049221:2046204],tree_1[2052239:2049222],tree_1[2055257:2052240],tree_2[1367153:1364136],tree_2[1370171:1367154]);
csa_3018 csau_3018_i730(tree_1[2058275:2055258],tree_1[2061293:2058276],tree_1[2064311:2061294],tree_2[1373189:1370172],tree_2[1376207:1373190]);
csa_3018 csau_3018_i731(tree_1[2067329:2064312],tree_1[2070347:2067330],tree_1[2073365:2070348],tree_2[1379225:1376208],tree_2[1382243:1379226]);
csa_3018 csau_3018_i732(tree_1[2076383:2073366],tree_1[2079401:2076384],tree_1[2082419:2079402],tree_2[1385261:1382244],tree_2[1388279:1385262]);
csa_3018 csau_3018_i733(tree_1[2085437:2082420],tree_1[2088455:2085438],tree_1[2091473:2088456],tree_2[1391297:1388280],tree_2[1394315:1391298]);
csa_3018 csau_3018_i734(tree_1[2094491:2091474],tree_1[2097509:2094492],tree_1[2100527:2097510],tree_2[1397333:1394316],tree_2[1400351:1397334]);
csa_3018 csau_3018_i735(tree_1[2103545:2100528],tree_1[2106563:2103546],tree_1[2109581:2106564],tree_2[1403369:1400352],tree_2[1406387:1403370]);
csa_3018 csau_3018_i736(tree_1[2112599:2109582],tree_1[2115617:2112600],tree_1[2118635:2115618],tree_2[1409405:1406388],tree_2[1412423:1409406]);
csa_3018 csau_3018_i737(tree_1[2121653:2118636],tree_1[2124671:2121654],tree_1[2127689:2124672],tree_2[1415441:1412424],tree_2[1418459:1415442]);
csa_3018 csau_3018_i738(tree_1[2130707:2127690],tree_1[2133725:2130708],tree_1[2136743:2133726],tree_2[1421477:1418460],tree_2[1424495:1421478]);
csa_3018 csau_3018_i739(tree_1[2139761:2136744],tree_1[2142779:2139762],tree_1[2145797:2142780],tree_2[1427513:1424496],tree_2[1430531:1427514]);
csa_3018 csau_3018_i740(tree_1[2148815:2145798],tree_1[2151833:2148816],tree_1[2154851:2151834],tree_2[1433549:1430532],tree_2[1436567:1433550]);
csa_3018 csau_3018_i741(tree_1[2157869:2154852],tree_1[2160887:2157870],tree_1[2163905:2160888],tree_2[1439585:1436568],tree_2[1442603:1439586]);
csa_3018 csau_3018_i742(tree_1[2166923:2163906],tree_1[2169941:2166924],tree_1[2172959:2169942],tree_2[1445621:1442604],tree_2[1448639:1445622]);
csa_3018 csau_3018_i743(tree_1[2175977:2172960],tree_1[2178995:2175978],tree_1[2182013:2178996],tree_2[1451657:1448640],tree_2[1454675:1451658]);
csa_3018 csau_3018_i744(tree_1[2185031:2182014],tree_1[2188049:2185032],tree_1[2191067:2188050],tree_2[1457693:1454676],tree_2[1460711:1457694]);
csa_3018 csau_3018_i745(tree_1[2194085:2191068],tree_1[2197103:2194086],tree_1[2200121:2197104],tree_2[1463729:1460712],tree_2[1466747:1463730]);
csa_3018 csau_3018_i746(tree_1[2203139:2200122],tree_1[2206157:2203140],tree_1[2209175:2206158],tree_2[1469765:1466748],tree_2[1472783:1469766]);
csa_3018 csau_3018_i747(tree_1[2212193:2209176],tree_1[2215211:2212194],tree_1[2218229:2215212],tree_2[1475801:1472784],tree_2[1478819:1475802]);
csa_3018 csau_3018_i748(tree_1[2221247:2218230],tree_1[2224265:2221248],tree_1[2227283:2224266],tree_2[1481837:1478820],tree_2[1484855:1481838]);
csa_3018 csau_3018_i749(tree_1[2230301:2227284],tree_1[2233319:2230302],tree_1[2236337:2233320],tree_2[1487873:1484856],tree_2[1490891:1487874]);
csa_3018 csau_3018_i750(tree_1[2239355:2236338],tree_1[2242373:2239356],tree_1[2245391:2242374],tree_2[1493909:1490892],tree_2[1496927:1493910]);
csa_3018 csau_3018_i751(tree_1[2248409:2245392],tree_1[2251427:2248410],tree_1[2254445:2251428],tree_2[1499945:1496928],tree_2[1502963:1499946]);
csa_3018 csau_3018_i752(tree_1[2257463:2254446],tree_1[2260481:2257464],tree_1[2263499:2260482],tree_2[1505981:1502964],tree_2[1508999:1505982]);
csa_3018 csau_3018_i753(tree_1[2266517:2263500],tree_1[2269535:2266518],tree_1[2272553:2269536],tree_2[1512017:1509000],tree_2[1515035:1512018]);
csa_3018 csau_3018_i754(tree_1[2275571:2272554],tree_1[2278589:2275572],tree_1[2281607:2278590],tree_2[1518053:1515036],tree_2[1521071:1518054]);
csa_3018 csau_3018_i755(tree_1[2284625:2281608],tree_1[2287643:2284626],tree_1[2290661:2287644],tree_2[1524089:1521072],tree_2[1527107:1524090]);
csa_3018 csau_3018_i756(tree_1[2293679:2290662],tree_1[2296697:2293680],tree_1[2299715:2296698],tree_2[1530125:1527108],tree_2[1533143:1530126]);
csa_3018 csau_3018_i757(tree_1[2302733:2299716],tree_1[2305751:2302734],tree_1[2308769:2305752],tree_2[1536161:1533144],tree_2[1539179:1536162]);
csa_3018 csau_3018_i758(tree_1[2311787:2308770],tree_1[2314805:2311788],tree_1[2317823:2314806],tree_2[1542197:1539180],tree_2[1545215:1542198]);
csa_3018 csau_3018_i759(tree_1[2320841:2317824],tree_1[2323859:2320842],tree_1[2326877:2323860],tree_2[1548233:1545216],tree_2[1551251:1548234]);
csa_3018 csau_3018_i760(tree_1[2329895:2326878],tree_1[2332913:2329896],tree_1[2335931:2332914],tree_2[1554269:1551252],tree_2[1557287:1554270]);
csa_3018 csau_3018_i761(tree_1[2338949:2335932],tree_1[2341967:2338950],tree_1[2344985:2341968],tree_2[1560305:1557288],tree_2[1563323:1560306]);
csa_3018 csau_3018_i762(tree_1[2348003:2344986],tree_1[2351021:2348004],tree_1[2354039:2351022],tree_2[1566341:1563324],tree_2[1569359:1566342]);
csa_3018 csau_3018_i763(tree_1[2357057:2354040],tree_1[2360075:2357058],tree_1[2363093:2360076],tree_2[1572377:1569360],tree_2[1575395:1572378]);
csa_3018 csau_3018_i764(tree_1[2366111:2363094],tree_1[2369129:2366112],tree_1[2372147:2369130],tree_2[1578413:1575396],tree_2[1581431:1578414]);
csa_3018 csau_3018_i765(tree_1[2375165:2372148],tree_1[2378183:2375166],tree_1[2381201:2378184],tree_2[1584449:1581432],tree_2[1587467:1584450]);
csa_3018 csau_3018_i766(tree_1[2384219:2381202],tree_1[2387237:2384220],tree_1[2390255:2387238],tree_2[1590485:1587468],tree_2[1593503:1590486]);
csa_3018 csau_3018_i767(tree_1[2393273:2390256],tree_1[2396291:2393274],tree_1[2399309:2396292],tree_2[1596521:1593504],tree_2[1599539:1596522]);
csa_3018 csau_3018_i768(tree_1[2402327:2399310],tree_1[2405345:2402328],tree_1[2408363:2405346],tree_2[1602557:1599540],tree_2[1605575:1602558]);
csa_3018 csau_3018_i769(tree_1[2411381:2408364],tree_1[2414399:2411382],tree_1[2417417:2414400],tree_2[1608593:1605576],tree_2[1611611:1608594]);
csa_3018 csau_3018_i770(tree_1[2420435:2417418],tree_1[2423453:2420436],tree_1[2426471:2423454],tree_2[1614629:1611612],tree_2[1617647:1614630]);
csa_3018 csau_3018_i771(tree_1[2429489:2426472],tree_1[2432507:2429490],tree_1[2435525:2432508],tree_2[1620665:1617648],tree_2[1623683:1620666]);
csa_3018 csau_3018_i772(tree_1[2438543:2435526],tree_1[2441561:2438544],tree_1[2444579:2441562],tree_2[1626701:1623684],tree_2[1629719:1626702]);
csa_3018 csau_3018_i773(tree_1[2447597:2444580],tree_1[2450615:2447598],tree_1[2453633:2450616],tree_2[1632737:1629720],tree_2[1635755:1632738]);
csa_3018 csau_3018_i774(tree_1[2456651:2453634],tree_1[2459669:2456652],tree_1[2462687:2459670],tree_2[1638773:1635756],tree_2[1641791:1638774]);
csa_3018 csau_3018_i775(tree_1[2465705:2462688],tree_1[2468723:2465706],tree_1[2471741:2468724],tree_2[1644809:1641792],tree_2[1647827:1644810]);
csa_3018 csau_3018_i776(tree_1[2474759:2471742],tree_1[2477777:2474760],tree_1[2480795:2477778],tree_2[1650845:1647828],tree_2[1653863:1650846]);
csa_3018 csau_3018_i777(tree_1[2483813:2480796],tree_1[2486831:2483814],tree_1[2489849:2486832],tree_2[1656881:1653864],tree_2[1659899:1656882]);
csa_3018 csau_3018_i778(tree_1[2492867:2489850],tree_1[2495885:2492868],tree_1[2498903:2495886],tree_2[1662917:1659900],tree_2[1665935:1662918]);
csa_3018 csau_3018_i779(tree_1[2501921:2498904],tree_1[2504939:2501922],tree_1[2507957:2504940],tree_2[1668953:1665936],tree_2[1671971:1668954]);
csa_3018 csau_3018_i780(tree_1[2510975:2507958],tree_1[2513993:2510976],tree_1[2517011:2513994],tree_2[1674989:1671972],tree_2[1678007:1674990]);
csa_3018 csau_3018_i781(tree_1[2520029:2517012],tree_1[2523047:2520030],tree_1[2526065:2523048],tree_2[1681025:1678008],tree_2[1684043:1681026]);
csa_3018 csau_3018_i782(tree_1[2529083:2526066],tree_1[2532101:2529084],tree_1[2535119:2532102],tree_2[1687061:1684044],tree_2[1690079:1687062]);
csa_3018 csau_3018_i783(tree_1[2538137:2535120],tree_1[2541155:2538138],tree_1[2544173:2541156],tree_2[1693097:1690080],tree_2[1696115:1693098]);
csa_3018 csau_3018_i784(tree_1[2547191:2544174],tree_1[2550209:2547192],tree_1[2553227:2550210],tree_2[1699133:1696116],tree_2[1702151:1699134]);
csa_3018 csau_3018_i785(tree_1[2556245:2553228],tree_1[2559263:2556246],tree_1[2562281:2559264],tree_2[1705169:1702152],tree_2[1708187:1705170]);
csa_3018 csau_3018_i786(tree_1[2565299:2562282],tree_1[2568317:2565300],tree_1[2571335:2568318],tree_2[1711205:1708188],tree_2[1714223:1711206]);
csa_3018 csau_3018_i787(tree_1[2574353:2571336],tree_1[2577371:2574354],tree_1[2580389:2577372],tree_2[1717241:1714224],tree_2[1720259:1717242]);
csa_3018 csau_3018_i788(tree_1[2583407:2580390],tree_1[2586425:2583408],tree_1[2589443:2586426],tree_2[1723277:1720260],tree_2[1726295:1723278]);
csa_3018 csau_3018_i789(tree_1[2592461:2589444],tree_1[2595479:2592462],tree_1[2598497:2595480],tree_2[1729313:1726296],tree_2[1732331:1729314]);
csa_3018 csau_3018_i790(tree_1[2601515:2598498],tree_1[2604533:2601516],tree_1[2607551:2604534],tree_2[1735349:1732332],tree_2[1738367:1735350]);
csa_3018 csau_3018_i791(tree_1[2610569:2607552],tree_1[2613587:2610570],tree_1[2616605:2613588],tree_2[1741385:1738368],tree_2[1744403:1741386]);
csa_3018 csau_3018_i792(tree_1[2619623:2616606],tree_1[2622641:2619624],tree_1[2625659:2622642],tree_2[1747421:1744404],tree_2[1750439:1747422]);
csa_3018 csau_3018_i793(tree_1[2628677:2625660],tree_1[2631695:2628678],tree_1[2634713:2631696],tree_2[1753457:1750440],tree_2[1756475:1753458]);
csa_3018 csau_3018_i794(tree_1[2637731:2634714],tree_1[2640749:2637732],tree_1[2643767:2640750],tree_2[1759493:1756476],tree_2[1762511:1759494]);
csa_3018 csau_3018_i795(tree_1[2646785:2643768],tree_1[2649803:2646786],tree_1[2652821:2649804],tree_2[1765529:1762512],tree_2[1768547:1765530]);
csa_3018 csau_3018_i796(tree_1[2655839:2652822],tree_1[2658857:2655840],tree_1[2661875:2658858],tree_2[1771565:1768548],tree_2[1774583:1771566]);
csa_3018 csau_3018_i797(tree_1[2664893:2661876],tree_1[2667911:2664894],tree_1[2670929:2667912],tree_2[1777601:1774584],tree_2[1780619:1777602]);
csa_3018 csau_3018_i798(tree_1[2673947:2670930],tree_1[2676965:2673948],tree_1[2679983:2676966],tree_2[1783637:1780620],tree_2[1786655:1783638]);
csa_3018 csau_3018_i799(tree_1[2683001:2679984],tree_1[2686019:2683002],tree_1[2689037:2686020],tree_2[1789673:1786656],tree_2[1792691:1789674]);
csa_3018 csau_3018_i800(tree_1[2692055:2689038],tree_1[2695073:2692056],tree_1[2698091:2695074],tree_2[1795709:1792692],tree_2[1798727:1795710]);
csa_3018 csau_3018_i801(tree_1[2701109:2698092],tree_1[2704127:2701110],tree_1[2707145:2704128],tree_2[1801745:1798728],tree_2[1804763:1801746]);
csa_3018 csau_3018_i802(tree_1[2710163:2707146],tree_1[2713181:2710164],tree_1[2716199:2713182],tree_2[1807781:1804764],tree_2[1810799:1807782]);
csa_3018 csau_3018_i803(tree_1[2719217:2716200],tree_1[2722235:2719218],tree_1[2725253:2722236],tree_2[1813817:1810800],tree_2[1816835:1813818]);
csa_3018 csau_3018_i804(tree_1[2728271:2725254],tree_1[2731289:2728272],tree_1[2734307:2731290],tree_2[1819853:1816836],tree_2[1822871:1819854]);
csa_3018 csau_3018_i805(tree_1[2737325:2734308],tree_1[2740343:2737326],tree_1[2743361:2740344],tree_2[1825889:1822872],tree_2[1828907:1825890]);
csa_3018 csau_3018_i806(tree_1[2746379:2743362],tree_1[2749397:2746380],tree_1[2752415:2749398],tree_2[1831925:1828908],tree_2[1834943:1831926]);
csa_3018 csau_3018_i807(tree_1[2755433:2752416],tree_1[2758451:2755434],tree_1[2761469:2758452],tree_2[1837961:1834944],tree_2[1840979:1837962]);
csa_3018 csau_3018_i808(tree_1[2764487:2761470],tree_1[2767505:2764488],tree_1[2770523:2767506],tree_2[1843997:1840980],tree_2[1847015:1843998]);
csa_3018 csau_3018_i809(tree_1[2773541:2770524],tree_1[2776559:2773542],tree_1[2779577:2776560],tree_2[1850033:1847016],tree_2[1853051:1850034]);
csa_3018 csau_3018_i810(tree_1[2782595:2779578],tree_1[2785613:2782596],tree_1[2788631:2785614],tree_2[1856069:1853052],tree_2[1859087:1856070]);
csa_3018 csau_3018_i811(tree_1[2791649:2788632],tree_1[2794667:2791650],tree_1[2797685:2794668],tree_2[1862105:1859088],tree_2[1865123:1862106]);
csa_3018 csau_3018_i812(tree_1[2800703:2797686],tree_1[2803721:2800704],tree_1[2806739:2803722],tree_2[1868141:1865124],tree_2[1871159:1868142]);
csa_3018 csau_3018_i813(tree_1[2809757:2806740],tree_1[2812775:2809758],tree_1[2815793:2812776],tree_2[1874177:1871160],tree_2[1877195:1874178]);
csa_3018 csau_3018_i814(tree_1[2818811:2815794],tree_1[2821829:2818812],tree_1[2824847:2821830],tree_2[1880213:1877196],tree_2[1883231:1880214]);
csa_3018 csau_3018_i815(tree_1[2827865:2824848],tree_1[2830883:2827866],tree_1[2833901:2830884],tree_2[1886249:1883232],tree_2[1889267:1886250]);
csa_3018 csau_3018_i816(tree_1[2836919:2833902],tree_1[2839937:2836920],tree_1[2842955:2839938],tree_2[1892285:1889268],tree_2[1895303:1892286]);
csa_3018 csau_3018_i817(tree_1[2845973:2842956],tree_1[2848991:2845974],tree_1[2852009:2848992],tree_2[1898321:1895304],tree_2[1901339:1898322]);
csa_3018 csau_3018_i818(tree_1[2855027:2852010],tree_1[2858045:2855028],tree_1[2861063:2858046],tree_2[1904357:1901340],tree_2[1907375:1904358]);
csa_3018 csau_3018_i819(tree_1[2864081:2861064],tree_1[2867099:2864082],tree_1[2870117:2867100],tree_2[1910393:1907376],tree_2[1913411:1910394]);
csa_3018 csau_3018_i820(tree_1[2873135:2870118],tree_1[2876153:2873136],tree_1[2879171:2876154],tree_2[1916429:1913412],tree_2[1919447:1916430]);
csa_3018 csau_3018_i821(tree_1[2882189:2879172],tree_1[2885207:2882190],tree_1[2888225:2885208],tree_2[1922465:1919448],tree_2[1925483:1922466]);
csa_3018 csau_3018_i822(tree_1[2891243:2888226],tree_1[2894261:2891244],tree_1[2897279:2894262],tree_2[1928501:1925484],tree_2[1931519:1928502]);
csa_3018 csau_3018_i823(tree_1[2900297:2897280],tree_1[2903315:2900298],tree_1[2906333:2903316],tree_2[1934537:1931520],tree_2[1937555:1934538]);
csa_3018 csau_3018_i824(tree_1[2909351:2906334],tree_1[2912369:2909352],tree_1[2915387:2912370],tree_2[1940573:1937556],tree_2[1943591:1940574]);
csa_3018 csau_3018_i825(tree_1[2918405:2915388],tree_1[2921423:2918406],tree_1[2924441:2921424],tree_2[1946609:1943592],tree_2[1949627:1946610]);
csa_3018 csau_3018_i826(tree_1[2927459:2924442],tree_1[2930477:2927460],tree_1[2933495:2930478],tree_2[1952645:1949628],tree_2[1955663:1952646]);
csa_3018 csau_3018_i827(tree_1[2936513:2933496],tree_1[2939531:2936514],tree_1[2942549:2939532],tree_2[1958681:1955664],tree_2[1961699:1958682]);
csa_3018 csau_3018_i828(tree_1[2945567:2942550],tree_1[2948585:2945568],tree_1[2951603:2948586],tree_2[1964717:1961700],tree_2[1967735:1964718]);
csa_3018 csau_3018_i829(tree_1[2954621:2951604],tree_1[2957639:2954622],tree_1[2960657:2957640],tree_2[1970753:1967736],tree_2[1973771:1970754]);
csa_3018 csau_3018_i830(tree_1[2963675:2960658],tree_1[2966693:2963676],tree_1[2969711:2966694],tree_2[1976789:1973772],tree_2[1979807:1976790]);
csa_3018 csau_3018_i831(tree_1[2972729:2969712],tree_1[2975747:2972730],tree_1[2978765:2975748],tree_2[1982825:1979808],tree_2[1985843:1982826]);
csa_3018 csau_3018_i832(tree_1[2981783:2978766],tree_1[2984801:2981784],tree_1[2987819:2984802],tree_2[1988861:1985844],tree_2[1991879:1988862]);
csa_3018 csau_3018_i833(tree_1[2990837:2987820],tree_1[2993855:2990838],tree_1[2996873:2993856],tree_2[1994897:1991880],tree_2[1997915:1994898]);
csa_3018 csau_3018_i834(tree_1[2999891:2996874],tree_1[3002909:2999892],tree_1[3005927:3002910],tree_2[2000933:1997916],tree_2[2003951:2000934]);
csa_3018 csau_3018_i835(tree_1[3008945:3005928],tree_1[3011963:3008946],tree_1[3014981:3011964],tree_2[2006969:2003952],tree_2[2009987:2006970]);
csa_3018 csau_3018_i836(tree_1[3017999:3014982],tree_1[3021017:3018000],tree_1[3024035:3021018],tree_2[2013005:2009988],tree_2[2016023:2013006]);
csa_3018 csau_3018_i837(tree_1[3027053:3024036],tree_1[3030071:3027054],tree_1[3033089:3030072],tree_2[2019041:2016024],tree_2[2022059:2019042]);
assign tree_2[2025077:2022060] = tree_1[3036107:3033090];
// layer-3
csa_3018 csau_3018_i838(tree_2[3017:0],tree_2[6035:3018],tree_2[9053:6036],tree_3[3017:0],tree_3[6035:3018]);
csa_3018 csau_3018_i839(tree_2[12071:9054],tree_2[15089:12072],tree_2[18107:15090],tree_3[9053:6036],tree_3[12071:9054]);
csa_3018 csau_3018_i840(tree_2[21125:18108],tree_2[24143:21126],tree_2[27161:24144],tree_3[15089:12072],tree_3[18107:15090]);
csa_3018 csau_3018_i841(tree_2[30179:27162],tree_2[33197:30180],tree_2[36215:33198],tree_3[21125:18108],tree_3[24143:21126]);
csa_3018 csau_3018_i842(tree_2[39233:36216],tree_2[42251:39234],tree_2[45269:42252],tree_3[27161:24144],tree_3[30179:27162]);
csa_3018 csau_3018_i843(tree_2[48287:45270],tree_2[51305:48288],tree_2[54323:51306],tree_3[33197:30180],tree_3[36215:33198]);
csa_3018 csau_3018_i844(tree_2[57341:54324],tree_2[60359:57342],tree_2[63377:60360],tree_3[39233:36216],tree_3[42251:39234]);
csa_3018 csau_3018_i845(tree_2[66395:63378],tree_2[69413:66396],tree_2[72431:69414],tree_3[45269:42252],tree_3[48287:45270]);
csa_3018 csau_3018_i846(tree_2[75449:72432],tree_2[78467:75450],tree_2[81485:78468],tree_3[51305:48288],tree_3[54323:51306]);
csa_3018 csau_3018_i847(tree_2[84503:81486],tree_2[87521:84504],tree_2[90539:87522],tree_3[57341:54324],tree_3[60359:57342]);
csa_3018 csau_3018_i848(tree_2[93557:90540],tree_2[96575:93558],tree_2[99593:96576],tree_3[63377:60360],tree_3[66395:63378]);
csa_3018 csau_3018_i849(tree_2[102611:99594],tree_2[105629:102612],tree_2[108647:105630],tree_3[69413:66396],tree_3[72431:69414]);
csa_3018 csau_3018_i850(tree_2[111665:108648],tree_2[114683:111666],tree_2[117701:114684],tree_3[75449:72432],tree_3[78467:75450]);
csa_3018 csau_3018_i851(tree_2[120719:117702],tree_2[123737:120720],tree_2[126755:123738],tree_3[81485:78468],tree_3[84503:81486]);
csa_3018 csau_3018_i852(tree_2[129773:126756],tree_2[132791:129774],tree_2[135809:132792],tree_3[87521:84504],tree_3[90539:87522]);
csa_3018 csau_3018_i853(tree_2[138827:135810],tree_2[141845:138828],tree_2[144863:141846],tree_3[93557:90540],tree_3[96575:93558]);
csa_3018 csau_3018_i854(tree_2[147881:144864],tree_2[150899:147882],tree_2[153917:150900],tree_3[99593:96576],tree_3[102611:99594]);
csa_3018 csau_3018_i855(tree_2[156935:153918],tree_2[159953:156936],tree_2[162971:159954],tree_3[105629:102612],tree_3[108647:105630]);
csa_3018 csau_3018_i856(tree_2[165989:162972],tree_2[169007:165990],tree_2[172025:169008],tree_3[111665:108648],tree_3[114683:111666]);
csa_3018 csau_3018_i857(tree_2[175043:172026],tree_2[178061:175044],tree_2[181079:178062],tree_3[117701:114684],tree_3[120719:117702]);
csa_3018 csau_3018_i858(tree_2[184097:181080],tree_2[187115:184098],tree_2[190133:187116],tree_3[123737:120720],tree_3[126755:123738]);
csa_3018 csau_3018_i859(tree_2[193151:190134],tree_2[196169:193152],tree_2[199187:196170],tree_3[129773:126756],tree_3[132791:129774]);
csa_3018 csau_3018_i860(tree_2[202205:199188],tree_2[205223:202206],tree_2[208241:205224],tree_3[135809:132792],tree_3[138827:135810]);
csa_3018 csau_3018_i861(tree_2[211259:208242],tree_2[214277:211260],tree_2[217295:214278],tree_3[141845:138828],tree_3[144863:141846]);
csa_3018 csau_3018_i862(tree_2[220313:217296],tree_2[223331:220314],tree_2[226349:223332],tree_3[147881:144864],tree_3[150899:147882]);
csa_3018 csau_3018_i863(tree_2[229367:226350],tree_2[232385:229368],tree_2[235403:232386],tree_3[153917:150900],tree_3[156935:153918]);
csa_3018 csau_3018_i864(tree_2[238421:235404],tree_2[241439:238422],tree_2[244457:241440],tree_3[159953:156936],tree_3[162971:159954]);
csa_3018 csau_3018_i865(tree_2[247475:244458],tree_2[250493:247476],tree_2[253511:250494],tree_3[165989:162972],tree_3[169007:165990]);
csa_3018 csau_3018_i866(tree_2[256529:253512],tree_2[259547:256530],tree_2[262565:259548],tree_3[172025:169008],tree_3[175043:172026]);
csa_3018 csau_3018_i867(tree_2[265583:262566],tree_2[268601:265584],tree_2[271619:268602],tree_3[178061:175044],tree_3[181079:178062]);
csa_3018 csau_3018_i868(tree_2[274637:271620],tree_2[277655:274638],tree_2[280673:277656],tree_3[184097:181080],tree_3[187115:184098]);
csa_3018 csau_3018_i869(tree_2[283691:280674],tree_2[286709:283692],tree_2[289727:286710],tree_3[190133:187116],tree_3[193151:190134]);
csa_3018 csau_3018_i870(tree_2[292745:289728],tree_2[295763:292746],tree_2[298781:295764],tree_3[196169:193152],tree_3[199187:196170]);
csa_3018 csau_3018_i871(tree_2[301799:298782],tree_2[304817:301800],tree_2[307835:304818],tree_3[202205:199188],tree_3[205223:202206]);
csa_3018 csau_3018_i872(tree_2[310853:307836],tree_2[313871:310854],tree_2[316889:313872],tree_3[208241:205224],tree_3[211259:208242]);
csa_3018 csau_3018_i873(tree_2[319907:316890],tree_2[322925:319908],tree_2[325943:322926],tree_3[214277:211260],tree_3[217295:214278]);
csa_3018 csau_3018_i874(tree_2[328961:325944],tree_2[331979:328962],tree_2[334997:331980],tree_3[220313:217296],tree_3[223331:220314]);
csa_3018 csau_3018_i875(tree_2[338015:334998],tree_2[341033:338016],tree_2[344051:341034],tree_3[226349:223332],tree_3[229367:226350]);
csa_3018 csau_3018_i876(tree_2[347069:344052],tree_2[350087:347070],tree_2[353105:350088],tree_3[232385:229368],tree_3[235403:232386]);
csa_3018 csau_3018_i877(tree_2[356123:353106],tree_2[359141:356124],tree_2[362159:359142],tree_3[238421:235404],tree_3[241439:238422]);
csa_3018 csau_3018_i878(tree_2[365177:362160],tree_2[368195:365178],tree_2[371213:368196],tree_3[244457:241440],tree_3[247475:244458]);
csa_3018 csau_3018_i879(tree_2[374231:371214],tree_2[377249:374232],tree_2[380267:377250],tree_3[250493:247476],tree_3[253511:250494]);
csa_3018 csau_3018_i880(tree_2[383285:380268],tree_2[386303:383286],tree_2[389321:386304],tree_3[256529:253512],tree_3[259547:256530]);
csa_3018 csau_3018_i881(tree_2[392339:389322],tree_2[395357:392340],tree_2[398375:395358],tree_3[262565:259548],tree_3[265583:262566]);
csa_3018 csau_3018_i882(tree_2[401393:398376],tree_2[404411:401394],tree_2[407429:404412],tree_3[268601:265584],tree_3[271619:268602]);
csa_3018 csau_3018_i883(tree_2[410447:407430],tree_2[413465:410448],tree_2[416483:413466],tree_3[274637:271620],tree_3[277655:274638]);
csa_3018 csau_3018_i884(tree_2[419501:416484],tree_2[422519:419502],tree_2[425537:422520],tree_3[280673:277656],tree_3[283691:280674]);
csa_3018 csau_3018_i885(tree_2[428555:425538],tree_2[431573:428556],tree_2[434591:431574],tree_3[286709:283692],tree_3[289727:286710]);
csa_3018 csau_3018_i886(tree_2[437609:434592],tree_2[440627:437610],tree_2[443645:440628],tree_3[292745:289728],tree_3[295763:292746]);
csa_3018 csau_3018_i887(tree_2[446663:443646],tree_2[449681:446664],tree_2[452699:449682],tree_3[298781:295764],tree_3[301799:298782]);
csa_3018 csau_3018_i888(tree_2[455717:452700],tree_2[458735:455718],tree_2[461753:458736],tree_3[304817:301800],tree_3[307835:304818]);
csa_3018 csau_3018_i889(tree_2[464771:461754],tree_2[467789:464772],tree_2[470807:467790],tree_3[310853:307836],tree_3[313871:310854]);
csa_3018 csau_3018_i890(tree_2[473825:470808],tree_2[476843:473826],tree_2[479861:476844],tree_3[316889:313872],tree_3[319907:316890]);
csa_3018 csau_3018_i891(tree_2[482879:479862],tree_2[485897:482880],tree_2[488915:485898],tree_3[322925:319908],tree_3[325943:322926]);
csa_3018 csau_3018_i892(tree_2[491933:488916],tree_2[494951:491934],tree_2[497969:494952],tree_3[328961:325944],tree_3[331979:328962]);
csa_3018 csau_3018_i893(tree_2[500987:497970],tree_2[504005:500988],tree_2[507023:504006],tree_3[334997:331980],tree_3[338015:334998]);
csa_3018 csau_3018_i894(tree_2[510041:507024],tree_2[513059:510042],tree_2[516077:513060],tree_3[341033:338016],tree_3[344051:341034]);
csa_3018 csau_3018_i895(tree_2[519095:516078],tree_2[522113:519096],tree_2[525131:522114],tree_3[347069:344052],tree_3[350087:347070]);
csa_3018 csau_3018_i896(tree_2[528149:525132],tree_2[531167:528150],tree_2[534185:531168],tree_3[353105:350088],tree_3[356123:353106]);
csa_3018 csau_3018_i897(tree_2[537203:534186],tree_2[540221:537204],tree_2[543239:540222],tree_3[359141:356124],tree_3[362159:359142]);
csa_3018 csau_3018_i898(tree_2[546257:543240],tree_2[549275:546258],tree_2[552293:549276],tree_3[365177:362160],tree_3[368195:365178]);
csa_3018 csau_3018_i899(tree_2[555311:552294],tree_2[558329:555312],tree_2[561347:558330],tree_3[371213:368196],tree_3[374231:371214]);
csa_3018 csau_3018_i900(tree_2[564365:561348],tree_2[567383:564366],tree_2[570401:567384],tree_3[377249:374232],tree_3[380267:377250]);
csa_3018 csau_3018_i901(tree_2[573419:570402],tree_2[576437:573420],tree_2[579455:576438],tree_3[383285:380268],tree_3[386303:383286]);
csa_3018 csau_3018_i902(tree_2[582473:579456],tree_2[585491:582474],tree_2[588509:585492],tree_3[389321:386304],tree_3[392339:389322]);
csa_3018 csau_3018_i903(tree_2[591527:588510],tree_2[594545:591528],tree_2[597563:594546],tree_3[395357:392340],tree_3[398375:395358]);
csa_3018 csau_3018_i904(tree_2[600581:597564],tree_2[603599:600582],tree_2[606617:603600],tree_3[401393:398376],tree_3[404411:401394]);
csa_3018 csau_3018_i905(tree_2[609635:606618],tree_2[612653:609636],tree_2[615671:612654],tree_3[407429:404412],tree_3[410447:407430]);
csa_3018 csau_3018_i906(tree_2[618689:615672],tree_2[621707:618690],tree_2[624725:621708],tree_3[413465:410448],tree_3[416483:413466]);
csa_3018 csau_3018_i907(tree_2[627743:624726],tree_2[630761:627744],tree_2[633779:630762],tree_3[419501:416484],tree_3[422519:419502]);
csa_3018 csau_3018_i908(tree_2[636797:633780],tree_2[639815:636798],tree_2[642833:639816],tree_3[425537:422520],tree_3[428555:425538]);
csa_3018 csau_3018_i909(tree_2[645851:642834],tree_2[648869:645852],tree_2[651887:648870],tree_3[431573:428556],tree_3[434591:431574]);
csa_3018 csau_3018_i910(tree_2[654905:651888],tree_2[657923:654906],tree_2[660941:657924],tree_3[437609:434592],tree_3[440627:437610]);
csa_3018 csau_3018_i911(tree_2[663959:660942],tree_2[666977:663960],tree_2[669995:666978],tree_3[443645:440628],tree_3[446663:443646]);
csa_3018 csau_3018_i912(tree_2[673013:669996],tree_2[676031:673014],tree_2[679049:676032],tree_3[449681:446664],tree_3[452699:449682]);
csa_3018 csau_3018_i913(tree_2[682067:679050],tree_2[685085:682068],tree_2[688103:685086],tree_3[455717:452700],tree_3[458735:455718]);
csa_3018 csau_3018_i914(tree_2[691121:688104],tree_2[694139:691122],tree_2[697157:694140],tree_3[461753:458736],tree_3[464771:461754]);
csa_3018 csau_3018_i915(tree_2[700175:697158],tree_2[703193:700176],tree_2[706211:703194],tree_3[467789:464772],tree_3[470807:467790]);
csa_3018 csau_3018_i916(tree_2[709229:706212],tree_2[712247:709230],tree_2[715265:712248],tree_3[473825:470808],tree_3[476843:473826]);
csa_3018 csau_3018_i917(tree_2[718283:715266],tree_2[721301:718284],tree_2[724319:721302],tree_3[479861:476844],tree_3[482879:479862]);
csa_3018 csau_3018_i918(tree_2[727337:724320],tree_2[730355:727338],tree_2[733373:730356],tree_3[485897:482880],tree_3[488915:485898]);
csa_3018 csau_3018_i919(tree_2[736391:733374],tree_2[739409:736392],tree_2[742427:739410],tree_3[491933:488916],tree_3[494951:491934]);
csa_3018 csau_3018_i920(tree_2[745445:742428],tree_2[748463:745446],tree_2[751481:748464],tree_3[497969:494952],tree_3[500987:497970]);
csa_3018 csau_3018_i921(tree_2[754499:751482],tree_2[757517:754500],tree_2[760535:757518],tree_3[504005:500988],tree_3[507023:504006]);
csa_3018 csau_3018_i922(tree_2[763553:760536],tree_2[766571:763554],tree_2[769589:766572],tree_3[510041:507024],tree_3[513059:510042]);
csa_3018 csau_3018_i923(tree_2[772607:769590],tree_2[775625:772608],tree_2[778643:775626],tree_3[516077:513060],tree_3[519095:516078]);
csa_3018 csau_3018_i924(tree_2[781661:778644],tree_2[784679:781662],tree_2[787697:784680],tree_3[522113:519096],tree_3[525131:522114]);
csa_3018 csau_3018_i925(tree_2[790715:787698],tree_2[793733:790716],tree_2[796751:793734],tree_3[528149:525132],tree_3[531167:528150]);
csa_3018 csau_3018_i926(tree_2[799769:796752],tree_2[802787:799770],tree_2[805805:802788],tree_3[534185:531168],tree_3[537203:534186]);
csa_3018 csau_3018_i927(tree_2[808823:805806],tree_2[811841:808824],tree_2[814859:811842],tree_3[540221:537204],tree_3[543239:540222]);
csa_3018 csau_3018_i928(tree_2[817877:814860],tree_2[820895:817878],tree_2[823913:820896],tree_3[546257:543240],tree_3[549275:546258]);
csa_3018 csau_3018_i929(tree_2[826931:823914],tree_2[829949:826932],tree_2[832967:829950],tree_3[552293:549276],tree_3[555311:552294]);
csa_3018 csau_3018_i930(tree_2[835985:832968],tree_2[839003:835986],tree_2[842021:839004],tree_3[558329:555312],tree_3[561347:558330]);
csa_3018 csau_3018_i931(tree_2[845039:842022],tree_2[848057:845040],tree_2[851075:848058],tree_3[564365:561348],tree_3[567383:564366]);
csa_3018 csau_3018_i932(tree_2[854093:851076],tree_2[857111:854094],tree_2[860129:857112],tree_3[570401:567384],tree_3[573419:570402]);
csa_3018 csau_3018_i933(tree_2[863147:860130],tree_2[866165:863148],tree_2[869183:866166],tree_3[576437:573420],tree_3[579455:576438]);
csa_3018 csau_3018_i934(tree_2[872201:869184],tree_2[875219:872202],tree_2[878237:875220],tree_3[582473:579456],tree_3[585491:582474]);
csa_3018 csau_3018_i935(tree_2[881255:878238],tree_2[884273:881256],tree_2[887291:884274],tree_3[588509:585492],tree_3[591527:588510]);
csa_3018 csau_3018_i936(tree_2[890309:887292],tree_2[893327:890310],tree_2[896345:893328],tree_3[594545:591528],tree_3[597563:594546]);
csa_3018 csau_3018_i937(tree_2[899363:896346],tree_2[902381:899364],tree_2[905399:902382],tree_3[600581:597564],tree_3[603599:600582]);
csa_3018 csau_3018_i938(tree_2[908417:905400],tree_2[911435:908418],tree_2[914453:911436],tree_3[606617:603600],tree_3[609635:606618]);
csa_3018 csau_3018_i939(tree_2[917471:914454],tree_2[920489:917472],tree_2[923507:920490],tree_3[612653:609636],tree_3[615671:612654]);
csa_3018 csau_3018_i940(tree_2[926525:923508],tree_2[929543:926526],tree_2[932561:929544],tree_3[618689:615672],tree_3[621707:618690]);
csa_3018 csau_3018_i941(tree_2[935579:932562],tree_2[938597:935580],tree_2[941615:938598],tree_3[624725:621708],tree_3[627743:624726]);
csa_3018 csau_3018_i942(tree_2[944633:941616],tree_2[947651:944634],tree_2[950669:947652],tree_3[630761:627744],tree_3[633779:630762]);
csa_3018 csau_3018_i943(tree_2[953687:950670],tree_2[956705:953688],tree_2[959723:956706],tree_3[636797:633780],tree_3[639815:636798]);
csa_3018 csau_3018_i944(tree_2[962741:959724],tree_2[965759:962742],tree_2[968777:965760],tree_3[642833:639816],tree_3[645851:642834]);
csa_3018 csau_3018_i945(tree_2[971795:968778],tree_2[974813:971796],tree_2[977831:974814],tree_3[648869:645852],tree_3[651887:648870]);
csa_3018 csau_3018_i946(tree_2[980849:977832],tree_2[983867:980850],tree_2[986885:983868],tree_3[654905:651888],tree_3[657923:654906]);
csa_3018 csau_3018_i947(tree_2[989903:986886],tree_2[992921:989904],tree_2[995939:992922],tree_3[660941:657924],tree_3[663959:660942]);
csa_3018 csau_3018_i948(tree_2[998957:995940],tree_2[1001975:998958],tree_2[1004993:1001976],tree_3[666977:663960],tree_3[669995:666978]);
csa_3018 csau_3018_i949(tree_2[1008011:1004994],tree_2[1011029:1008012],tree_2[1014047:1011030],tree_3[673013:669996],tree_3[676031:673014]);
csa_3018 csau_3018_i950(tree_2[1017065:1014048],tree_2[1020083:1017066],tree_2[1023101:1020084],tree_3[679049:676032],tree_3[682067:679050]);
csa_3018 csau_3018_i951(tree_2[1026119:1023102],tree_2[1029137:1026120],tree_2[1032155:1029138],tree_3[685085:682068],tree_3[688103:685086]);
csa_3018 csau_3018_i952(tree_2[1035173:1032156],tree_2[1038191:1035174],tree_2[1041209:1038192],tree_3[691121:688104],tree_3[694139:691122]);
csa_3018 csau_3018_i953(tree_2[1044227:1041210],tree_2[1047245:1044228],tree_2[1050263:1047246],tree_3[697157:694140],tree_3[700175:697158]);
csa_3018 csau_3018_i954(tree_2[1053281:1050264],tree_2[1056299:1053282],tree_2[1059317:1056300],tree_3[703193:700176],tree_3[706211:703194]);
csa_3018 csau_3018_i955(tree_2[1062335:1059318],tree_2[1065353:1062336],tree_2[1068371:1065354],tree_3[709229:706212],tree_3[712247:709230]);
csa_3018 csau_3018_i956(tree_2[1071389:1068372],tree_2[1074407:1071390],tree_2[1077425:1074408],tree_3[715265:712248],tree_3[718283:715266]);
csa_3018 csau_3018_i957(tree_2[1080443:1077426],tree_2[1083461:1080444],tree_2[1086479:1083462],tree_3[721301:718284],tree_3[724319:721302]);
csa_3018 csau_3018_i958(tree_2[1089497:1086480],tree_2[1092515:1089498],tree_2[1095533:1092516],tree_3[727337:724320],tree_3[730355:727338]);
csa_3018 csau_3018_i959(tree_2[1098551:1095534],tree_2[1101569:1098552],tree_2[1104587:1101570],tree_3[733373:730356],tree_3[736391:733374]);
csa_3018 csau_3018_i960(tree_2[1107605:1104588],tree_2[1110623:1107606],tree_2[1113641:1110624],tree_3[739409:736392],tree_3[742427:739410]);
csa_3018 csau_3018_i961(tree_2[1116659:1113642],tree_2[1119677:1116660],tree_2[1122695:1119678],tree_3[745445:742428],tree_3[748463:745446]);
csa_3018 csau_3018_i962(tree_2[1125713:1122696],tree_2[1128731:1125714],tree_2[1131749:1128732],tree_3[751481:748464],tree_3[754499:751482]);
csa_3018 csau_3018_i963(tree_2[1134767:1131750],tree_2[1137785:1134768],tree_2[1140803:1137786],tree_3[757517:754500],tree_3[760535:757518]);
csa_3018 csau_3018_i964(tree_2[1143821:1140804],tree_2[1146839:1143822],tree_2[1149857:1146840],tree_3[763553:760536],tree_3[766571:763554]);
csa_3018 csau_3018_i965(tree_2[1152875:1149858],tree_2[1155893:1152876],tree_2[1158911:1155894],tree_3[769589:766572],tree_3[772607:769590]);
csa_3018 csau_3018_i966(tree_2[1161929:1158912],tree_2[1164947:1161930],tree_2[1167965:1164948],tree_3[775625:772608],tree_3[778643:775626]);
csa_3018 csau_3018_i967(tree_2[1170983:1167966],tree_2[1174001:1170984],tree_2[1177019:1174002],tree_3[781661:778644],tree_3[784679:781662]);
csa_3018 csau_3018_i968(tree_2[1180037:1177020],tree_2[1183055:1180038],tree_2[1186073:1183056],tree_3[787697:784680],tree_3[790715:787698]);
csa_3018 csau_3018_i969(tree_2[1189091:1186074],tree_2[1192109:1189092],tree_2[1195127:1192110],tree_3[793733:790716],tree_3[796751:793734]);
csa_3018 csau_3018_i970(tree_2[1198145:1195128],tree_2[1201163:1198146],tree_2[1204181:1201164],tree_3[799769:796752],tree_3[802787:799770]);
csa_3018 csau_3018_i971(tree_2[1207199:1204182],tree_2[1210217:1207200],tree_2[1213235:1210218],tree_3[805805:802788],tree_3[808823:805806]);
csa_3018 csau_3018_i972(tree_2[1216253:1213236],tree_2[1219271:1216254],tree_2[1222289:1219272],tree_3[811841:808824],tree_3[814859:811842]);
csa_3018 csau_3018_i973(tree_2[1225307:1222290],tree_2[1228325:1225308],tree_2[1231343:1228326],tree_3[817877:814860],tree_3[820895:817878]);
csa_3018 csau_3018_i974(tree_2[1234361:1231344],tree_2[1237379:1234362],tree_2[1240397:1237380],tree_3[823913:820896],tree_3[826931:823914]);
csa_3018 csau_3018_i975(tree_2[1243415:1240398],tree_2[1246433:1243416],tree_2[1249451:1246434],tree_3[829949:826932],tree_3[832967:829950]);
csa_3018 csau_3018_i976(tree_2[1252469:1249452],tree_2[1255487:1252470],tree_2[1258505:1255488],tree_3[835985:832968],tree_3[839003:835986]);
csa_3018 csau_3018_i977(tree_2[1261523:1258506],tree_2[1264541:1261524],tree_2[1267559:1264542],tree_3[842021:839004],tree_3[845039:842022]);
csa_3018 csau_3018_i978(tree_2[1270577:1267560],tree_2[1273595:1270578],tree_2[1276613:1273596],tree_3[848057:845040],tree_3[851075:848058]);
csa_3018 csau_3018_i979(tree_2[1279631:1276614],tree_2[1282649:1279632],tree_2[1285667:1282650],tree_3[854093:851076],tree_3[857111:854094]);
csa_3018 csau_3018_i980(tree_2[1288685:1285668],tree_2[1291703:1288686],tree_2[1294721:1291704],tree_3[860129:857112],tree_3[863147:860130]);
csa_3018 csau_3018_i981(tree_2[1297739:1294722],tree_2[1300757:1297740],tree_2[1303775:1300758],tree_3[866165:863148],tree_3[869183:866166]);
csa_3018 csau_3018_i982(tree_2[1306793:1303776],tree_2[1309811:1306794],tree_2[1312829:1309812],tree_3[872201:869184],tree_3[875219:872202]);
csa_3018 csau_3018_i983(tree_2[1315847:1312830],tree_2[1318865:1315848],tree_2[1321883:1318866],tree_3[878237:875220],tree_3[881255:878238]);
csa_3018 csau_3018_i984(tree_2[1324901:1321884],tree_2[1327919:1324902],tree_2[1330937:1327920],tree_3[884273:881256],tree_3[887291:884274]);
csa_3018 csau_3018_i985(tree_2[1333955:1330938],tree_2[1336973:1333956],tree_2[1339991:1336974],tree_3[890309:887292],tree_3[893327:890310]);
csa_3018 csau_3018_i986(tree_2[1343009:1339992],tree_2[1346027:1343010],tree_2[1349045:1346028],tree_3[896345:893328],tree_3[899363:896346]);
csa_3018 csau_3018_i987(tree_2[1352063:1349046],tree_2[1355081:1352064],tree_2[1358099:1355082],tree_3[902381:899364],tree_3[905399:902382]);
csa_3018 csau_3018_i988(tree_2[1361117:1358100],tree_2[1364135:1361118],tree_2[1367153:1364136],tree_3[908417:905400],tree_3[911435:908418]);
csa_3018 csau_3018_i989(tree_2[1370171:1367154],tree_2[1373189:1370172],tree_2[1376207:1373190],tree_3[914453:911436],tree_3[917471:914454]);
csa_3018 csau_3018_i990(tree_2[1379225:1376208],tree_2[1382243:1379226],tree_2[1385261:1382244],tree_3[920489:917472],tree_3[923507:920490]);
csa_3018 csau_3018_i991(tree_2[1388279:1385262],tree_2[1391297:1388280],tree_2[1394315:1391298],tree_3[926525:923508],tree_3[929543:926526]);
csa_3018 csau_3018_i992(tree_2[1397333:1394316],tree_2[1400351:1397334],tree_2[1403369:1400352],tree_3[932561:929544],tree_3[935579:932562]);
csa_3018 csau_3018_i993(tree_2[1406387:1403370],tree_2[1409405:1406388],tree_2[1412423:1409406],tree_3[938597:935580],tree_3[941615:938598]);
csa_3018 csau_3018_i994(tree_2[1415441:1412424],tree_2[1418459:1415442],tree_2[1421477:1418460],tree_3[944633:941616],tree_3[947651:944634]);
csa_3018 csau_3018_i995(tree_2[1424495:1421478],tree_2[1427513:1424496],tree_2[1430531:1427514],tree_3[950669:947652],tree_3[953687:950670]);
csa_3018 csau_3018_i996(tree_2[1433549:1430532],tree_2[1436567:1433550],tree_2[1439585:1436568],tree_3[956705:953688],tree_3[959723:956706]);
csa_3018 csau_3018_i997(tree_2[1442603:1439586],tree_2[1445621:1442604],tree_2[1448639:1445622],tree_3[962741:959724],tree_3[965759:962742]);
csa_3018 csau_3018_i998(tree_2[1451657:1448640],tree_2[1454675:1451658],tree_2[1457693:1454676],tree_3[968777:965760],tree_3[971795:968778]);
csa_3018 csau_3018_i999(tree_2[1460711:1457694],tree_2[1463729:1460712],tree_2[1466747:1463730],tree_3[974813:971796],tree_3[977831:974814]);
csa_3018 csau_3018_i1000(tree_2[1469765:1466748],tree_2[1472783:1469766],tree_2[1475801:1472784],tree_3[980849:977832],tree_3[983867:980850]);
csa_3018 csau_3018_i1001(tree_2[1478819:1475802],tree_2[1481837:1478820],tree_2[1484855:1481838],tree_3[986885:983868],tree_3[989903:986886]);
csa_3018 csau_3018_i1002(tree_2[1487873:1484856],tree_2[1490891:1487874],tree_2[1493909:1490892],tree_3[992921:989904],tree_3[995939:992922]);
csa_3018 csau_3018_i1003(tree_2[1496927:1493910],tree_2[1499945:1496928],tree_2[1502963:1499946],tree_3[998957:995940],tree_3[1001975:998958]);
csa_3018 csau_3018_i1004(tree_2[1505981:1502964],tree_2[1508999:1505982],tree_2[1512017:1509000],tree_3[1004993:1001976],tree_3[1008011:1004994]);
csa_3018 csau_3018_i1005(tree_2[1515035:1512018],tree_2[1518053:1515036],tree_2[1521071:1518054],tree_3[1011029:1008012],tree_3[1014047:1011030]);
csa_3018 csau_3018_i1006(tree_2[1524089:1521072],tree_2[1527107:1524090],tree_2[1530125:1527108],tree_3[1017065:1014048],tree_3[1020083:1017066]);
csa_3018 csau_3018_i1007(tree_2[1533143:1530126],tree_2[1536161:1533144],tree_2[1539179:1536162],tree_3[1023101:1020084],tree_3[1026119:1023102]);
csa_3018 csau_3018_i1008(tree_2[1542197:1539180],tree_2[1545215:1542198],tree_2[1548233:1545216],tree_3[1029137:1026120],tree_3[1032155:1029138]);
csa_3018 csau_3018_i1009(tree_2[1551251:1548234],tree_2[1554269:1551252],tree_2[1557287:1554270],tree_3[1035173:1032156],tree_3[1038191:1035174]);
csa_3018 csau_3018_i1010(tree_2[1560305:1557288],tree_2[1563323:1560306],tree_2[1566341:1563324],tree_3[1041209:1038192],tree_3[1044227:1041210]);
csa_3018 csau_3018_i1011(tree_2[1569359:1566342],tree_2[1572377:1569360],tree_2[1575395:1572378],tree_3[1047245:1044228],tree_3[1050263:1047246]);
csa_3018 csau_3018_i1012(tree_2[1578413:1575396],tree_2[1581431:1578414],tree_2[1584449:1581432],tree_3[1053281:1050264],tree_3[1056299:1053282]);
csa_3018 csau_3018_i1013(tree_2[1587467:1584450],tree_2[1590485:1587468],tree_2[1593503:1590486],tree_3[1059317:1056300],tree_3[1062335:1059318]);
csa_3018 csau_3018_i1014(tree_2[1596521:1593504],tree_2[1599539:1596522],tree_2[1602557:1599540],tree_3[1065353:1062336],tree_3[1068371:1065354]);
csa_3018 csau_3018_i1015(tree_2[1605575:1602558],tree_2[1608593:1605576],tree_2[1611611:1608594],tree_3[1071389:1068372],tree_3[1074407:1071390]);
csa_3018 csau_3018_i1016(tree_2[1614629:1611612],tree_2[1617647:1614630],tree_2[1620665:1617648],tree_3[1077425:1074408],tree_3[1080443:1077426]);
csa_3018 csau_3018_i1017(tree_2[1623683:1620666],tree_2[1626701:1623684],tree_2[1629719:1626702],tree_3[1083461:1080444],tree_3[1086479:1083462]);
csa_3018 csau_3018_i1018(tree_2[1632737:1629720],tree_2[1635755:1632738],tree_2[1638773:1635756],tree_3[1089497:1086480],tree_3[1092515:1089498]);
csa_3018 csau_3018_i1019(tree_2[1641791:1638774],tree_2[1644809:1641792],tree_2[1647827:1644810],tree_3[1095533:1092516],tree_3[1098551:1095534]);
csa_3018 csau_3018_i1020(tree_2[1650845:1647828],tree_2[1653863:1650846],tree_2[1656881:1653864],tree_3[1101569:1098552],tree_3[1104587:1101570]);
csa_3018 csau_3018_i1021(tree_2[1659899:1656882],tree_2[1662917:1659900],tree_2[1665935:1662918],tree_3[1107605:1104588],tree_3[1110623:1107606]);
csa_3018 csau_3018_i1022(tree_2[1668953:1665936],tree_2[1671971:1668954],tree_2[1674989:1671972],tree_3[1113641:1110624],tree_3[1116659:1113642]);
csa_3018 csau_3018_i1023(tree_2[1678007:1674990],tree_2[1681025:1678008],tree_2[1684043:1681026],tree_3[1119677:1116660],tree_3[1122695:1119678]);
csa_3018 csau_3018_i1024(tree_2[1687061:1684044],tree_2[1690079:1687062],tree_2[1693097:1690080],tree_3[1125713:1122696],tree_3[1128731:1125714]);
csa_3018 csau_3018_i1025(tree_2[1696115:1693098],tree_2[1699133:1696116],tree_2[1702151:1699134],tree_3[1131749:1128732],tree_3[1134767:1131750]);
csa_3018 csau_3018_i1026(tree_2[1705169:1702152],tree_2[1708187:1705170],tree_2[1711205:1708188],tree_3[1137785:1134768],tree_3[1140803:1137786]);
csa_3018 csau_3018_i1027(tree_2[1714223:1711206],tree_2[1717241:1714224],tree_2[1720259:1717242],tree_3[1143821:1140804],tree_3[1146839:1143822]);
csa_3018 csau_3018_i1028(tree_2[1723277:1720260],tree_2[1726295:1723278],tree_2[1729313:1726296],tree_3[1149857:1146840],tree_3[1152875:1149858]);
csa_3018 csau_3018_i1029(tree_2[1732331:1729314],tree_2[1735349:1732332],tree_2[1738367:1735350],tree_3[1155893:1152876],tree_3[1158911:1155894]);
csa_3018 csau_3018_i1030(tree_2[1741385:1738368],tree_2[1744403:1741386],tree_2[1747421:1744404],tree_3[1161929:1158912],tree_3[1164947:1161930]);
csa_3018 csau_3018_i1031(tree_2[1750439:1747422],tree_2[1753457:1750440],tree_2[1756475:1753458],tree_3[1167965:1164948],tree_3[1170983:1167966]);
csa_3018 csau_3018_i1032(tree_2[1759493:1756476],tree_2[1762511:1759494],tree_2[1765529:1762512],tree_3[1174001:1170984],tree_3[1177019:1174002]);
csa_3018 csau_3018_i1033(tree_2[1768547:1765530],tree_2[1771565:1768548],tree_2[1774583:1771566],tree_3[1180037:1177020],tree_3[1183055:1180038]);
csa_3018 csau_3018_i1034(tree_2[1777601:1774584],tree_2[1780619:1777602],tree_2[1783637:1780620],tree_3[1186073:1183056],tree_3[1189091:1186074]);
csa_3018 csau_3018_i1035(tree_2[1786655:1783638],tree_2[1789673:1786656],tree_2[1792691:1789674],tree_3[1192109:1189092],tree_3[1195127:1192110]);
csa_3018 csau_3018_i1036(tree_2[1795709:1792692],tree_2[1798727:1795710],tree_2[1801745:1798728],tree_3[1198145:1195128],tree_3[1201163:1198146]);
csa_3018 csau_3018_i1037(tree_2[1804763:1801746],tree_2[1807781:1804764],tree_2[1810799:1807782],tree_3[1204181:1201164],tree_3[1207199:1204182]);
csa_3018 csau_3018_i1038(tree_2[1813817:1810800],tree_2[1816835:1813818],tree_2[1819853:1816836],tree_3[1210217:1207200],tree_3[1213235:1210218]);
csa_3018 csau_3018_i1039(tree_2[1822871:1819854],tree_2[1825889:1822872],tree_2[1828907:1825890],tree_3[1216253:1213236],tree_3[1219271:1216254]);
csa_3018 csau_3018_i1040(tree_2[1831925:1828908],tree_2[1834943:1831926],tree_2[1837961:1834944],tree_3[1222289:1219272],tree_3[1225307:1222290]);
csa_3018 csau_3018_i1041(tree_2[1840979:1837962],tree_2[1843997:1840980],tree_2[1847015:1843998],tree_3[1228325:1225308],tree_3[1231343:1228326]);
csa_3018 csau_3018_i1042(tree_2[1850033:1847016],tree_2[1853051:1850034],tree_2[1856069:1853052],tree_3[1234361:1231344],tree_3[1237379:1234362]);
csa_3018 csau_3018_i1043(tree_2[1859087:1856070],tree_2[1862105:1859088],tree_2[1865123:1862106],tree_3[1240397:1237380],tree_3[1243415:1240398]);
csa_3018 csau_3018_i1044(tree_2[1868141:1865124],tree_2[1871159:1868142],tree_2[1874177:1871160],tree_3[1246433:1243416],tree_3[1249451:1246434]);
csa_3018 csau_3018_i1045(tree_2[1877195:1874178],tree_2[1880213:1877196],tree_2[1883231:1880214],tree_3[1252469:1249452],tree_3[1255487:1252470]);
csa_3018 csau_3018_i1046(tree_2[1886249:1883232],tree_2[1889267:1886250],tree_2[1892285:1889268],tree_3[1258505:1255488],tree_3[1261523:1258506]);
csa_3018 csau_3018_i1047(tree_2[1895303:1892286],tree_2[1898321:1895304],tree_2[1901339:1898322],tree_3[1264541:1261524],tree_3[1267559:1264542]);
csa_3018 csau_3018_i1048(tree_2[1904357:1901340],tree_2[1907375:1904358],tree_2[1910393:1907376],tree_3[1270577:1267560],tree_3[1273595:1270578]);
csa_3018 csau_3018_i1049(tree_2[1913411:1910394],tree_2[1916429:1913412],tree_2[1919447:1916430],tree_3[1276613:1273596],tree_3[1279631:1276614]);
csa_3018 csau_3018_i1050(tree_2[1922465:1919448],tree_2[1925483:1922466],tree_2[1928501:1925484],tree_3[1282649:1279632],tree_3[1285667:1282650]);
csa_3018 csau_3018_i1051(tree_2[1931519:1928502],tree_2[1934537:1931520],tree_2[1937555:1934538],tree_3[1288685:1285668],tree_3[1291703:1288686]);
csa_3018 csau_3018_i1052(tree_2[1940573:1937556],tree_2[1943591:1940574],tree_2[1946609:1943592],tree_3[1294721:1291704],tree_3[1297739:1294722]);
csa_3018 csau_3018_i1053(tree_2[1949627:1946610],tree_2[1952645:1949628],tree_2[1955663:1952646],tree_3[1300757:1297740],tree_3[1303775:1300758]);
csa_3018 csau_3018_i1054(tree_2[1958681:1955664],tree_2[1961699:1958682],tree_2[1964717:1961700],tree_3[1306793:1303776],tree_3[1309811:1306794]);
csa_3018 csau_3018_i1055(tree_2[1967735:1964718],tree_2[1970753:1967736],tree_2[1973771:1970754],tree_3[1312829:1309812],tree_3[1315847:1312830]);
csa_3018 csau_3018_i1056(tree_2[1976789:1973772],tree_2[1979807:1976790],tree_2[1982825:1979808],tree_3[1318865:1315848],tree_3[1321883:1318866]);
csa_3018 csau_3018_i1057(tree_2[1985843:1982826],tree_2[1988861:1985844],tree_2[1991879:1988862],tree_3[1324901:1321884],tree_3[1327919:1324902]);
csa_3018 csau_3018_i1058(tree_2[1994897:1991880],tree_2[1997915:1994898],tree_2[2000933:1997916],tree_3[1330937:1327920],tree_3[1333955:1330938]);
csa_3018 csau_3018_i1059(tree_2[2003951:2000934],tree_2[2006969:2003952],tree_2[2009987:2006970],tree_3[1336973:1333956],tree_3[1339991:1336974]);
csa_3018 csau_3018_i1060(tree_2[2013005:2009988],tree_2[2016023:2013006],tree_2[2019041:2016024],tree_3[1343009:1339992],tree_3[1346027:1343010]);
assign tree_3[1349045:1346028] = tree_2[2022059:2019042];
assign tree_3[1352063:1349046] = tree_2[2025077:2022060];
// layer-4
csa_3018 csau_3018_i1061(tree_3[3017:0],tree_3[6035:3018],tree_3[9053:6036],tree_4[3017:0],tree_4[6035:3018]);
csa_3018 csau_3018_i1062(tree_3[12071:9054],tree_3[15089:12072],tree_3[18107:15090],tree_4[9053:6036],tree_4[12071:9054]);
csa_3018 csau_3018_i1063(tree_3[21125:18108],tree_3[24143:21126],tree_3[27161:24144],tree_4[15089:12072],tree_4[18107:15090]);
csa_3018 csau_3018_i1064(tree_3[30179:27162],tree_3[33197:30180],tree_3[36215:33198],tree_4[21125:18108],tree_4[24143:21126]);
csa_3018 csau_3018_i1065(tree_3[39233:36216],tree_3[42251:39234],tree_3[45269:42252],tree_4[27161:24144],tree_4[30179:27162]);
csa_3018 csau_3018_i1066(tree_3[48287:45270],tree_3[51305:48288],tree_3[54323:51306],tree_4[33197:30180],tree_4[36215:33198]);
csa_3018 csau_3018_i1067(tree_3[57341:54324],tree_3[60359:57342],tree_3[63377:60360],tree_4[39233:36216],tree_4[42251:39234]);
csa_3018 csau_3018_i1068(tree_3[66395:63378],tree_3[69413:66396],tree_3[72431:69414],tree_4[45269:42252],tree_4[48287:45270]);
csa_3018 csau_3018_i1069(tree_3[75449:72432],tree_3[78467:75450],tree_3[81485:78468],tree_4[51305:48288],tree_4[54323:51306]);
csa_3018 csau_3018_i1070(tree_3[84503:81486],tree_3[87521:84504],tree_3[90539:87522],tree_4[57341:54324],tree_4[60359:57342]);
csa_3018 csau_3018_i1071(tree_3[93557:90540],tree_3[96575:93558],tree_3[99593:96576],tree_4[63377:60360],tree_4[66395:63378]);
csa_3018 csau_3018_i1072(tree_3[102611:99594],tree_3[105629:102612],tree_3[108647:105630],tree_4[69413:66396],tree_4[72431:69414]);
csa_3018 csau_3018_i1073(tree_3[111665:108648],tree_3[114683:111666],tree_3[117701:114684],tree_4[75449:72432],tree_4[78467:75450]);
csa_3018 csau_3018_i1074(tree_3[120719:117702],tree_3[123737:120720],tree_3[126755:123738],tree_4[81485:78468],tree_4[84503:81486]);
csa_3018 csau_3018_i1075(tree_3[129773:126756],tree_3[132791:129774],tree_3[135809:132792],tree_4[87521:84504],tree_4[90539:87522]);
csa_3018 csau_3018_i1076(tree_3[138827:135810],tree_3[141845:138828],tree_3[144863:141846],tree_4[93557:90540],tree_4[96575:93558]);
csa_3018 csau_3018_i1077(tree_3[147881:144864],tree_3[150899:147882],tree_3[153917:150900],tree_4[99593:96576],tree_4[102611:99594]);
csa_3018 csau_3018_i1078(tree_3[156935:153918],tree_3[159953:156936],tree_3[162971:159954],tree_4[105629:102612],tree_4[108647:105630]);
csa_3018 csau_3018_i1079(tree_3[165989:162972],tree_3[169007:165990],tree_3[172025:169008],tree_4[111665:108648],tree_4[114683:111666]);
csa_3018 csau_3018_i1080(tree_3[175043:172026],tree_3[178061:175044],tree_3[181079:178062],tree_4[117701:114684],tree_4[120719:117702]);
csa_3018 csau_3018_i1081(tree_3[184097:181080],tree_3[187115:184098],tree_3[190133:187116],tree_4[123737:120720],tree_4[126755:123738]);
csa_3018 csau_3018_i1082(tree_3[193151:190134],tree_3[196169:193152],tree_3[199187:196170],tree_4[129773:126756],tree_4[132791:129774]);
csa_3018 csau_3018_i1083(tree_3[202205:199188],tree_3[205223:202206],tree_3[208241:205224],tree_4[135809:132792],tree_4[138827:135810]);
csa_3018 csau_3018_i1084(tree_3[211259:208242],tree_3[214277:211260],tree_3[217295:214278],tree_4[141845:138828],tree_4[144863:141846]);
csa_3018 csau_3018_i1085(tree_3[220313:217296],tree_3[223331:220314],tree_3[226349:223332],tree_4[147881:144864],tree_4[150899:147882]);
csa_3018 csau_3018_i1086(tree_3[229367:226350],tree_3[232385:229368],tree_3[235403:232386],tree_4[153917:150900],tree_4[156935:153918]);
csa_3018 csau_3018_i1087(tree_3[238421:235404],tree_3[241439:238422],tree_3[244457:241440],tree_4[159953:156936],tree_4[162971:159954]);
csa_3018 csau_3018_i1088(tree_3[247475:244458],tree_3[250493:247476],tree_3[253511:250494],tree_4[165989:162972],tree_4[169007:165990]);
csa_3018 csau_3018_i1089(tree_3[256529:253512],tree_3[259547:256530],tree_3[262565:259548],tree_4[172025:169008],tree_4[175043:172026]);
csa_3018 csau_3018_i1090(tree_3[265583:262566],tree_3[268601:265584],tree_3[271619:268602],tree_4[178061:175044],tree_4[181079:178062]);
csa_3018 csau_3018_i1091(tree_3[274637:271620],tree_3[277655:274638],tree_3[280673:277656],tree_4[184097:181080],tree_4[187115:184098]);
csa_3018 csau_3018_i1092(tree_3[283691:280674],tree_3[286709:283692],tree_3[289727:286710],tree_4[190133:187116],tree_4[193151:190134]);
csa_3018 csau_3018_i1093(tree_3[292745:289728],tree_3[295763:292746],tree_3[298781:295764],tree_4[196169:193152],tree_4[199187:196170]);
csa_3018 csau_3018_i1094(tree_3[301799:298782],tree_3[304817:301800],tree_3[307835:304818],tree_4[202205:199188],tree_4[205223:202206]);
csa_3018 csau_3018_i1095(tree_3[310853:307836],tree_3[313871:310854],tree_3[316889:313872],tree_4[208241:205224],tree_4[211259:208242]);
csa_3018 csau_3018_i1096(tree_3[319907:316890],tree_3[322925:319908],tree_3[325943:322926],tree_4[214277:211260],tree_4[217295:214278]);
csa_3018 csau_3018_i1097(tree_3[328961:325944],tree_3[331979:328962],tree_3[334997:331980],tree_4[220313:217296],tree_4[223331:220314]);
csa_3018 csau_3018_i1098(tree_3[338015:334998],tree_3[341033:338016],tree_3[344051:341034],tree_4[226349:223332],tree_4[229367:226350]);
csa_3018 csau_3018_i1099(tree_3[347069:344052],tree_3[350087:347070],tree_3[353105:350088],tree_4[232385:229368],tree_4[235403:232386]);
csa_3018 csau_3018_i1100(tree_3[356123:353106],tree_3[359141:356124],tree_3[362159:359142],tree_4[238421:235404],tree_4[241439:238422]);
csa_3018 csau_3018_i1101(tree_3[365177:362160],tree_3[368195:365178],tree_3[371213:368196],tree_4[244457:241440],tree_4[247475:244458]);
csa_3018 csau_3018_i1102(tree_3[374231:371214],tree_3[377249:374232],tree_3[380267:377250],tree_4[250493:247476],tree_4[253511:250494]);
csa_3018 csau_3018_i1103(tree_3[383285:380268],tree_3[386303:383286],tree_3[389321:386304],tree_4[256529:253512],tree_4[259547:256530]);
csa_3018 csau_3018_i1104(tree_3[392339:389322],tree_3[395357:392340],tree_3[398375:395358],tree_4[262565:259548],tree_4[265583:262566]);
csa_3018 csau_3018_i1105(tree_3[401393:398376],tree_3[404411:401394],tree_3[407429:404412],tree_4[268601:265584],tree_4[271619:268602]);
csa_3018 csau_3018_i1106(tree_3[410447:407430],tree_3[413465:410448],tree_3[416483:413466],tree_4[274637:271620],tree_4[277655:274638]);
csa_3018 csau_3018_i1107(tree_3[419501:416484],tree_3[422519:419502],tree_3[425537:422520],tree_4[280673:277656],tree_4[283691:280674]);
csa_3018 csau_3018_i1108(tree_3[428555:425538],tree_3[431573:428556],tree_3[434591:431574],tree_4[286709:283692],tree_4[289727:286710]);
csa_3018 csau_3018_i1109(tree_3[437609:434592],tree_3[440627:437610],tree_3[443645:440628],tree_4[292745:289728],tree_4[295763:292746]);
csa_3018 csau_3018_i1110(tree_3[446663:443646],tree_3[449681:446664],tree_3[452699:449682],tree_4[298781:295764],tree_4[301799:298782]);
csa_3018 csau_3018_i1111(tree_3[455717:452700],tree_3[458735:455718],tree_3[461753:458736],tree_4[304817:301800],tree_4[307835:304818]);
csa_3018 csau_3018_i1112(tree_3[464771:461754],tree_3[467789:464772],tree_3[470807:467790],tree_4[310853:307836],tree_4[313871:310854]);
csa_3018 csau_3018_i1113(tree_3[473825:470808],tree_3[476843:473826],tree_3[479861:476844],tree_4[316889:313872],tree_4[319907:316890]);
csa_3018 csau_3018_i1114(tree_3[482879:479862],tree_3[485897:482880],tree_3[488915:485898],tree_4[322925:319908],tree_4[325943:322926]);
csa_3018 csau_3018_i1115(tree_3[491933:488916],tree_3[494951:491934],tree_3[497969:494952],tree_4[328961:325944],tree_4[331979:328962]);
csa_3018 csau_3018_i1116(tree_3[500987:497970],tree_3[504005:500988],tree_3[507023:504006],tree_4[334997:331980],tree_4[338015:334998]);
csa_3018 csau_3018_i1117(tree_3[510041:507024],tree_3[513059:510042],tree_3[516077:513060],tree_4[341033:338016],tree_4[344051:341034]);
csa_3018 csau_3018_i1118(tree_3[519095:516078],tree_3[522113:519096],tree_3[525131:522114],tree_4[347069:344052],tree_4[350087:347070]);
csa_3018 csau_3018_i1119(tree_3[528149:525132],tree_3[531167:528150],tree_3[534185:531168],tree_4[353105:350088],tree_4[356123:353106]);
csa_3018 csau_3018_i1120(tree_3[537203:534186],tree_3[540221:537204],tree_3[543239:540222],tree_4[359141:356124],tree_4[362159:359142]);
csa_3018 csau_3018_i1121(tree_3[546257:543240],tree_3[549275:546258],tree_3[552293:549276],tree_4[365177:362160],tree_4[368195:365178]);
csa_3018 csau_3018_i1122(tree_3[555311:552294],tree_3[558329:555312],tree_3[561347:558330],tree_4[371213:368196],tree_4[374231:371214]);
csa_3018 csau_3018_i1123(tree_3[564365:561348],tree_3[567383:564366],tree_3[570401:567384],tree_4[377249:374232],tree_4[380267:377250]);
csa_3018 csau_3018_i1124(tree_3[573419:570402],tree_3[576437:573420],tree_3[579455:576438],tree_4[383285:380268],tree_4[386303:383286]);
csa_3018 csau_3018_i1125(tree_3[582473:579456],tree_3[585491:582474],tree_3[588509:585492],tree_4[389321:386304],tree_4[392339:389322]);
csa_3018 csau_3018_i1126(tree_3[591527:588510],tree_3[594545:591528],tree_3[597563:594546],tree_4[395357:392340],tree_4[398375:395358]);
csa_3018 csau_3018_i1127(tree_3[600581:597564],tree_3[603599:600582],tree_3[606617:603600],tree_4[401393:398376],tree_4[404411:401394]);
csa_3018 csau_3018_i1128(tree_3[609635:606618],tree_3[612653:609636],tree_3[615671:612654],tree_4[407429:404412],tree_4[410447:407430]);
csa_3018 csau_3018_i1129(tree_3[618689:615672],tree_3[621707:618690],tree_3[624725:621708],tree_4[413465:410448],tree_4[416483:413466]);
csa_3018 csau_3018_i1130(tree_3[627743:624726],tree_3[630761:627744],tree_3[633779:630762],tree_4[419501:416484],tree_4[422519:419502]);
csa_3018 csau_3018_i1131(tree_3[636797:633780],tree_3[639815:636798],tree_3[642833:639816],tree_4[425537:422520],tree_4[428555:425538]);
csa_3018 csau_3018_i1132(tree_3[645851:642834],tree_3[648869:645852],tree_3[651887:648870],tree_4[431573:428556],tree_4[434591:431574]);
csa_3018 csau_3018_i1133(tree_3[654905:651888],tree_3[657923:654906],tree_3[660941:657924],tree_4[437609:434592],tree_4[440627:437610]);
csa_3018 csau_3018_i1134(tree_3[663959:660942],tree_3[666977:663960],tree_3[669995:666978],tree_4[443645:440628],tree_4[446663:443646]);
csa_3018 csau_3018_i1135(tree_3[673013:669996],tree_3[676031:673014],tree_3[679049:676032],tree_4[449681:446664],tree_4[452699:449682]);
csa_3018 csau_3018_i1136(tree_3[682067:679050],tree_3[685085:682068],tree_3[688103:685086],tree_4[455717:452700],tree_4[458735:455718]);
csa_3018 csau_3018_i1137(tree_3[691121:688104],tree_3[694139:691122],tree_3[697157:694140],tree_4[461753:458736],tree_4[464771:461754]);
csa_3018 csau_3018_i1138(tree_3[700175:697158],tree_3[703193:700176],tree_3[706211:703194],tree_4[467789:464772],tree_4[470807:467790]);
csa_3018 csau_3018_i1139(tree_3[709229:706212],tree_3[712247:709230],tree_3[715265:712248],tree_4[473825:470808],tree_4[476843:473826]);
csa_3018 csau_3018_i1140(tree_3[718283:715266],tree_3[721301:718284],tree_3[724319:721302],tree_4[479861:476844],tree_4[482879:479862]);
csa_3018 csau_3018_i1141(tree_3[727337:724320],tree_3[730355:727338],tree_3[733373:730356],tree_4[485897:482880],tree_4[488915:485898]);
csa_3018 csau_3018_i1142(tree_3[736391:733374],tree_3[739409:736392],tree_3[742427:739410],tree_4[491933:488916],tree_4[494951:491934]);
csa_3018 csau_3018_i1143(tree_3[745445:742428],tree_3[748463:745446],tree_3[751481:748464],tree_4[497969:494952],tree_4[500987:497970]);
csa_3018 csau_3018_i1144(tree_3[754499:751482],tree_3[757517:754500],tree_3[760535:757518],tree_4[504005:500988],tree_4[507023:504006]);
csa_3018 csau_3018_i1145(tree_3[763553:760536],tree_3[766571:763554],tree_3[769589:766572],tree_4[510041:507024],tree_4[513059:510042]);
csa_3018 csau_3018_i1146(tree_3[772607:769590],tree_3[775625:772608],tree_3[778643:775626],tree_4[516077:513060],tree_4[519095:516078]);
csa_3018 csau_3018_i1147(tree_3[781661:778644],tree_3[784679:781662],tree_3[787697:784680],tree_4[522113:519096],tree_4[525131:522114]);
csa_3018 csau_3018_i1148(tree_3[790715:787698],tree_3[793733:790716],tree_3[796751:793734],tree_4[528149:525132],tree_4[531167:528150]);
csa_3018 csau_3018_i1149(tree_3[799769:796752],tree_3[802787:799770],tree_3[805805:802788],tree_4[534185:531168],tree_4[537203:534186]);
csa_3018 csau_3018_i1150(tree_3[808823:805806],tree_3[811841:808824],tree_3[814859:811842],tree_4[540221:537204],tree_4[543239:540222]);
csa_3018 csau_3018_i1151(tree_3[817877:814860],tree_3[820895:817878],tree_3[823913:820896],tree_4[546257:543240],tree_4[549275:546258]);
csa_3018 csau_3018_i1152(tree_3[826931:823914],tree_3[829949:826932],tree_3[832967:829950],tree_4[552293:549276],tree_4[555311:552294]);
csa_3018 csau_3018_i1153(tree_3[835985:832968],tree_3[839003:835986],tree_3[842021:839004],tree_4[558329:555312],tree_4[561347:558330]);
csa_3018 csau_3018_i1154(tree_3[845039:842022],tree_3[848057:845040],tree_3[851075:848058],tree_4[564365:561348],tree_4[567383:564366]);
csa_3018 csau_3018_i1155(tree_3[854093:851076],tree_3[857111:854094],tree_3[860129:857112],tree_4[570401:567384],tree_4[573419:570402]);
csa_3018 csau_3018_i1156(tree_3[863147:860130],tree_3[866165:863148],tree_3[869183:866166],tree_4[576437:573420],tree_4[579455:576438]);
csa_3018 csau_3018_i1157(tree_3[872201:869184],tree_3[875219:872202],tree_3[878237:875220],tree_4[582473:579456],tree_4[585491:582474]);
csa_3018 csau_3018_i1158(tree_3[881255:878238],tree_3[884273:881256],tree_3[887291:884274],tree_4[588509:585492],tree_4[591527:588510]);
csa_3018 csau_3018_i1159(tree_3[890309:887292],tree_3[893327:890310],tree_3[896345:893328],tree_4[594545:591528],tree_4[597563:594546]);
csa_3018 csau_3018_i1160(tree_3[899363:896346],tree_3[902381:899364],tree_3[905399:902382],tree_4[600581:597564],tree_4[603599:600582]);
csa_3018 csau_3018_i1161(tree_3[908417:905400],tree_3[911435:908418],tree_3[914453:911436],tree_4[606617:603600],tree_4[609635:606618]);
csa_3018 csau_3018_i1162(tree_3[917471:914454],tree_3[920489:917472],tree_3[923507:920490],tree_4[612653:609636],tree_4[615671:612654]);
csa_3018 csau_3018_i1163(tree_3[926525:923508],tree_3[929543:926526],tree_3[932561:929544],tree_4[618689:615672],tree_4[621707:618690]);
csa_3018 csau_3018_i1164(tree_3[935579:932562],tree_3[938597:935580],tree_3[941615:938598],tree_4[624725:621708],tree_4[627743:624726]);
csa_3018 csau_3018_i1165(tree_3[944633:941616],tree_3[947651:944634],tree_3[950669:947652],tree_4[630761:627744],tree_4[633779:630762]);
csa_3018 csau_3018_i1166(tree_3[953687:950670],tree_3[956705:953688],tree_3[959723:956706],tree_4[636797:633780],tree_4[639815:636798]);
csa_3018 csau_3018_i1167(tree_3[962741:959724],tree_3[965759:962742],tree_3[968777:965760],tree_4[642833:639816],tree_4[645851:642834]);
csa_3018 csau_3018_i1168(tree_3[971795:968778],tree_3[974813:971796],tree_3[977831:974814],tree_4[648869:645852],tree_4[651887:648870]);
csa_3018 csau_3018_i1169(tree_3[980849:977832],tree_3[983867:980850],tree_3[986885:983868],tree_4[654905:651888],tree_4[657923:654906]);
csa_3018 csau_3018_i1170(tree_3[989903:986886],tree_3[992921:989904],tree_3[995939:992922],tree_4[660941:657924],tree_4[663959:660942]);
csa_3018 csau_3018_i1171(tree_3[998957:995940],tree_3[1001975:998958],tree_3[1004993:1001976],tree_4[666977:663960],tree_4[669995:666978]);
csa_3018 csau_3018_i1172(tree_3[1008011:1004994],tree_3[1011029:1008012],tree_3[1014047:1011030],tree_4[673013:669996],tree_4[676031:673014]);
csa_3018 csau_3018_i1173(tree_3[1017065:1014048],tree_3[1020083:1017066],tree_3[1023101:1020084],tree_4[679049:676032],tree_4[682067:679050]);
csa_3018 csau_3018_i1174(tree_3[1026119:1023102],tree_3[1029137:1026120],tree_3[1032155:1029138],tree_4[685085:682068],tree_4[688103:685086]);
csa_3018 csau_3018_i1175(tree_3[1035173:1032156],tree_3[1038191:1035174],tree_3[1041209:1038192],tree_4[691121:688104],tree_4[694139:691122]);
csa_3018 csau_3018_i1176(tree_3[1044227:1041210],tree_3[1047245:1044228],tree_3[1050263:1047246],tree_4[697157:694140],tree_4[700175:697158]);
csa_3018 csau_3018_i1177(tree_3[1053281:1050264],tree_3[1056299:1053282],tree_3[1059317:1056300],tree_4[703193:700176],tree_4[706211:703194]);
csa_3018 csau_3018_i1178(tree_3[1062335:1059318],tree_3[1065353:1062336],tree_3[1068371:1065354],tree_4[709229:706212],tree_4[712247:709230]);
csa_3018 csau_3018_i1179(tree_3[1071389:1068372],tree_3[1074407:1071390],tree_3[1077425:1074408],tree_4[715265:712248],tree_4[718283:715266]);
csa_3018 csau_3018_i1180(tree_3[1080443:1077426],tree_3[1083461:1080444],tree_3[1086479:1083462],tree_4[721301:718284],tree_4[724319:721302]);
csa_3018 csau_3018_i1181(tree_3[1089497:1086480],tree_3[1092515:1089498],tree_3[1095533:1092516],tree_4[727337:724320],tree_4[730355:727338]);
csa_3018 csau_3018_i1182(tree_3[1098551:1095534],tree_3[1101569:1098552],tree_3[1104587:1101570],tree_4[733373:730356],tree_4[736391:733374]);
csa_3018 csau_3018_i1183(tree_3[1107605:1104588],tree_3[1110623:1107606],tree_3[1113641:1110624],tree_4[739409:736392],tree_4[742427:739410]);
csa_3018 csau_3018_i1184(tree_3[1116659:1113642],tree_3[1119677:1116660],tree_3[1122695:1119678],tree_4[745445:742428],tree_4[748463:745446]);
csa_3018 csau_3018_i1185(tree_3[1125713:1122696],tree_3[1128731:1125714],tree_3[1131749:1128732],tree_4[751481:748464],tree_4[754499:751482]);
csa_3018 csau_3018_i1186(tree_3[1134767:1131750],tree_3[1137785:1134768],tree_3[1140803:1137786],tree_4[757517:754500],tree_4[760535:757518]);
csa_3018 csau_3018_i1187(tree_3[1143821:1140804],tree_3[1146839:1143822],tree_3[1149857:1146840],tree_4[763553:760536],tree_4[766571:763554]);
csa_3018 csau_3018_i1188(tree_3[1152875:1149858],tree_3[1155893:1152876],tree_3[1158911:1155894],tree_4[769589:766572],tree_4[772607:769590]);
csa_3018 csau_3018_i1189(tree_3[1161929:1158912],tree_3[1164947:1161930],tree_3[1167965:1164948],tree_4[775625:772608],tree_4[778643:775626]);
csa_3018 csau_3018_i1190(tree_3[1170983:1167966],tree_3[1174001:1170984],tree_3[1177019:1174002],tree_4[781661:778644],tree_4[784679:781662]);
csa_3018 csau_3018_i1191(tree_3[1180037:1177020],tree_3[1183055:1180038],tree_3[1186073:1183056],tree_4[787697:784680],tree_4[790715:787698]);
csa_3018 csau_3018_i1192(tree_3[1189091:1186074],tree_3[1192109:1189092],tree_3[1195127:1192110],tree_4[793733:790716],tree_4[796751:793734]);
csa_3018 csau_3018_i1193(tree_3[1198145:1195128],tree_3[1201163:1198146],tree_3[1204181:1201164],tree_4[799769:796752],tree_4[802787:799770]);
csa_3018 csau_3018_i1194(tree_3[1207199:1204182],tree_3[1210217:1207200],tree_3[1213235:1210218],tree_4[805805:802788],tree_4[808823:805806]);
csa_3018 csau_3018_i1195(tree_3[1216253:1213236],tree_3[1219271:1216254],tree_3[1222289:1219272],tree_4[811841:808824],tree_4[814859:811842]);
csa_3018 csau_3018_i1196(tree_3[1225307:1222290],tree_3[1228325:1225308],tree_3[1231343:1228326],tree_4[817877:814860],tree_4[820895:817878]);
csa_3018 csau_3018_i1197(tree_3[1234361:1231344],tree_3[1237379:1234362],tree_3[1240397:1237380],tree_4[823913:820896],tree_4[826931:823914]);
csa_3018 csau_3018_i1198(tree_3[1243415:1240398],tree_3[1246433:1243416],tree_3[1249451:1246434],tree_4[829949:826932],tree_4[832967:829950]);
csa_3018 csau_3018_i1199(tree_3[1252469:1249452],tree_3[1255487:1252470],tree_3[1258505:1255488],tree_4[835985:832968],tree_4[839003:835986]);
csa_3018 csau_3018_i1200(tree_3[1261523:1258506],tree_3[1264541:1261524],tree_3[1267559:1264542],tree_4[842021:839004],tree_4[845039:842022]);
csa_3018 csau_3018_i1201(tree_3[1270577:1267560],tree_3[1273595:1270578],tree_3[1276613:1273596],tree_4[848057:845040],tree_4[851075:848058]);
csa_3018 csau_3018_i1202(tree_3[1279631:1276614],tree_3[1282649:1279632],tree_3[1285667:1282650],tree_4[854093:851076],tree_4[857111:854094]);
csa_3018 csau_3018_i1203(tree_3[1288685:1285668],tree_3[1291703:1288686],tree_3[1294721:1291704],tree_4[860129:857112],tree_4[863147:860130]);
csa_3018 csau_3018_i1204(tree_3[1297739:1294722],tree_3[1300757:1297740],tree_3[1303775:1300758],tree_4[866165:863148],tree_4[869183:866166]);
csa_3018 csau_3018_i1205(tree_3[1306793:1303776],tree_3[1309811:1306794],tree_3[1312829:1309812],tree_4[872201:869184],tree_4[875219:872202]);
csa_3018 csau_3018_i1206(tree_3[1315847:1312830],tree_3[1318865:1315848],tree_3[1321883:1318866],tree_4[878237:875220],tree_4[881255:878238]);
csa_3018 csau_3018_i1207(tree_3[1324901:1321884],tree_3[1327919:1324902],tree_3[1330937:1327920],tree_4[884273:881256],tree_4[887291:884274]);
csa_3018 csau_3018_i1208(tree_3[1333955:1330938],tree_3[1336973:1333956],tree_3[1339991:1336974],tree_4[890309:887292],tree_4[893327:890310]);
csa_3018 csau_3018_i1209(tree_3[1343009:1339992],tree_3[1346027:1343010],tree_3[1349045:1346028],tree_4[896345:893328],tree_4[899363:896346]);
assign tree_4[902381:899364] = tree_3[1352063:1349046];
// layer-5
csa_3018 csau_3018_i1210(tree_4[3017:0],tree_4[6035:3018],tree_4[9053:6036],tree_5[3017:0],tree_5[6035:3018]);
csa_3018 csau_3018_i1211(tree_4[12071:9054],tree_4[15089:12072],tree_4[18107:15090],tree_5[9053:6036],tree_5[12071:9054]);
csa_3018 csau_3018_i1212(tree_4[21125:18108],tree_4[24143:21126],tree_4[27161:24144],tree_5[15089:12072],tree_5[18107:15090]);
csa_3018 csau_3018_i1213(tree_4[30179:27162],tree_4[33197:30180],tree_4[36215:33198],tree_5[21125:18108],tree_5[24143:21126]);
csa_3018 csau_3018_i1214(tree_4[39233:36216],tree_4[42251:39234],tree_4[45269:42252],tree_5[27161:24144],tree_5[30179:27162]);
csa_3018 csau_3018_i1215(tree_4[48287:45270],tree_4[51305:48288],tree_4[54323:51306],tree_5[33197:30180],tree_5[36215:33198]);
csa_3018 csau_3018_i1216(tree_4[57341:54324],tree_4[60359:57342],tree_4[63377:60360],tree_5[39233:36216],tree_5[42251:39234]);
csa_3018 csau_3018_i1217(tree_4[66395:63378],tree_4[69413:66396],tree_4[72431:69414],tree_5[45269:42252],tree_5[48287:45270]);
csa_3018 csau_3018_i1218(tree_4[75449:72432],tree_4[78467:75450],tree_4[81485:78468],tree_5[51305:48288],tree_5[54323:51306]);
csa_3018 csau_3018_i1219(tree_4[84503:81486],tree_4[87521:84504],tree_4[90539:87522],tree_5[57341:54324],tree_5[60359:57342]);
csa_3018 csau_3018_i1220(tree_4[93557:90540],tree_4[96575:93558],tree_4[99593:96576],tree_5[63377:60360],tree_5[66395:63378]);
csa_3018 csau_3018_i1221(tree_4[102611:99594],tree_4[105629:102612],tree_4[108647:105630],tree_5[69413:66396],tree_5[72431:69414]);
csa_3018 csau_3018_i1222(tree_4[111665:108648],tree_4[114683:111666],tree_4[117701:114684],tree_5[75449:72432],tree_5[78467:75450]);
csa_3018 csau_3018_i1223(tree_4[120719:117702],tree_4[123737:120720],tree_4[126755:123738],tree_5[81485:78468],tree_5[84503:81486]);
csa_3018 csau_3018_i1224(tree_4[129773:126756],tree_4[132791:129774],tree_4[135809:132792],tree_5[87521:84504],tree_5[90539:87522]);
csa_3018 csau_3018_i1225(tree_4[138827:135810],tree_4[141845:138828],tree_4[144863:141846],tree_5[93557:90540],tree_5[96575:93558]);
csa_3018 csau_3018_i1226(tree_4[147881:144864],tree_4[150899:147882],tree_4[153917:150900],tree_5[99593:96576],tree_5[102611:99594]);
csa_3018 csau_3018_i1227(tree_4[156935:153918],tree_4[159953:156936],tree_4[162971:159954],tree_5[105629:102612],tree_5[108647:105630]);
csa_3018 csau_3018_i1228(tree_4[165989:162972],tree_4[169007:165990],tree_4[172025:169008],tree_5[111665:108648],tree_5[114683:111666]);
csa_3018 csau_3018_i1229(tree_4[175043:172026],tree_4[178061:175044],tree_4[181079:178062],tree_5[117701:114684],tree_5[120719:117702]);
csa_3018 csau_3018_i1230(tree_4[184097:181080],tree_4[187115:184098],tree_4[190133:187116],tree_5[123737:120720],tree_5[126755:123738]);
csa_3018 csau_3018_i1231(tree_4[193151:190134],tree_4[196169:193152],tree_4[199187:196170],tree_5[129773:126756],tree_5[132791:129774]);
csa_3018 csau_3018_i1232(tree_4[202205:199188],tree_4[205223:202206],tree_4[208241:205224],tree_5[135809:132792],tree_5[138827:135810]);
csa_3018 csau_3018_i1233(tree_4[211259:208242],tree_4[214277:211260],tree_4[217295:214278],tree_5[141845:138828],tree_5[144863:141846]);
csa_3018 csau_3018_i1234(tree_4[220313:217296],tree_4[223331:220314],tree_4[226349:223332],tree_5[147881:144864],tree_5[150899:147882]);
csa_3018 csau_3018_i1235(tree_4[229367:226350],tree_4[232385:229368],tree_4[235403:232386],tree_5[153917:150900],tree_5[156935:153918]);
csa_3018 csau_3018_i1236(tree_4[238421:235404],tree_4[241439:238422],tree_4[244457:241440],tree_5[159953:156936],tree_5[162971:159954]);
csa_3018 csau_3018_i1237(tree_4[247475:244458],tree_4[250493:247476],tree_4[253511:250494],tree_5[165989:162972],tree_5[169007:165990]);
csa_3018 csau_3018_i1238(tree_4[256529:253512],tree_4[259547:256530],tree_4[262565:259548],tree_5[172025:169008],tree_5[175043:172026]);
csa_3018 csau_3018_i1239(tree_4[265583:262566],tree_4[268601:265584],tree_4[271619:268602],tree_5[178061:175044],tree_5[181079:178062]);
csa_3018 csau_3018_i1240(tree_4[274637:271620],tree_4[277655:274638],tree_4[280673:277656],tree_5[184097:181080],tree_5[187115:184098]);
csa_3018 csau_3018_i1241(tree_4[283691:280674],tree_4[286709:283692],tree_4[289727:286710],tree_5[190133:187116],tree_5[193151:190134]);
csa_3018 csau_3018_i1242(tree_4[292745:289728],tree_4[295763:292746],tree_4[298781:295764],tree_5[196169:193152],tree_5[199187:196170]);
csa_3018 csau_3018_i1243(tree_4[301799:298782],tree_4[304817:301800],tree_4[307835:304818],tree_5[202205:199188],tree_5[205223:202206]);
csa_3018 csau_3018_i1244(tree_4[310853:307836],tree_4[313871:310854],tree_4[316889:313872],tree_5[208241:205224],tree_5[211259:208242]);
csa_3018 csau_3018_i1245(tree_4[319907:316890],tree_4[322925:319908],tree_4[325943:322926],tree_5[214277:211260],tree_5[217295:214278]);
csa_3018 csau_3018_i1246(tree_4[328961:325944],tree_4[331979:328962],tree_4[334997:331980],tree_5[220313:217296],tree_5[223331:220314]);
csa_3018 csau_3018_i1247(tree_4[338015:334998],tree_4[341033:338016],tree_4[344051:341034],tree_5[226349:223332],tree_5[229367:226350]);
csa_3018 csau_3018_i1248(tree_4[347069:344052],tree_4[350087:347070],tree_4[353105:350088],tree_5[232385:229368],tree_5[235403:232386]);
csa_3018 csau_3018_i1249(tree_4[356123:353106],tree_4[359141:356124],tree_4[362159:359142],tree_5[238421:235404],tree_5[241439:238422]);
csa_3018 csau_3018_i1250(tree_4[365177:362160],tree_4[368195:365178],tree_4[371213:368196],tree_5[244457:241440],tree_5[247475:244458]);
csa_3018 csau_3018_i1251(tree_4[374231:371214],tree_4[377249:374232],tree_4[380267:377250],tree_5[250493:247476],tree_5[253511:250494]);
csa_3018 csau_3018_i1252(tree_4[383285:380268],tree_4[386303:383286],tree_4[389321:386304],tree_5[256529:253512],tree_5[259547:256530]);
csa_3018 csau_3018_i1253(tree_4[392339:389322],tree_4[395357:392340],tree_4[398375:395358],tree_5[262565:259548],tree_5[265583:262566]);
csa_3018 csau_3018_i1254(tree_4[401393:398376],tree_4[404411:401394],tree_4[407429:404412],tree_5[268601:265584],tree_5[271619:268602]);
csa_3018 csau_3018_i1255(tree_4[410447:407430],tree_4[413465:410448],tree_4[416483:413466],tree_5[274637:271620],tree_5[277655:274638]);
csa_3018 csau_3018_i1256(tree_4[419501:416484],tree_4[422519:419502],tree_4[425537:422520],tree_5[280673:277656],tree_5[283691:280674]);
csa_3018 csau_3018_i1257(tree_4[428555:425538],tree_4[431573:428556],tree_4[434591:431574],tree_5[286709:283692],tree_5[289727:286710]);
csa_3018 csau_3018_i1258(tree_4[437609:434592],tree_4[440627:437610],tree_4[443645:440628],tree_5[292745:289728],tree_5[295763:292746]);
csa_3018 csau_3018_i1259(tree_4[446663:443646],tree_4[449681:446664],tree_4[452699:449682],tree_5[298781:295764],tree_5[301799:298782]);
csa_3018 csau_3018_i1260(tree_4[455717:452700],tree_4[458735:455718],tree_4[461753:458736],tree_5[304817:301800],tree_5[307835:304818]);
csa_3018 csau_3018_i1261(tree_4[464771:461754],tree_4[467789:464772],tree_4[470807:467790],tree_5[310853:307836],tree_5[313871:310854]);
csa_3018 csau_3018_i1262(tree_4[473825:470808],tree_4[476843:473826],tree_4[479861:476844],tree_5[316889:313872],tree_5[319907:316890]);
csa_3018 csau_3018_i1263(tree_4[482879:479862],tree_4[485897:482880],tree_4[488915:485898],tree_5[322925:319908],tree_5[325943:322926]);
csa_3018 csau_3018_i1264(tree_4[491933:488916],tree_4[494951:491934],tree_4[497969:494952],tree_5[328961:325944],tree_5[331979:328962]);
csa_3018 csau_3018_i1265(tree_4[500987:497970],tree_4[504005:500988],tree_4[507023:504006],tree_5[334997:331980],tree_5[338015:334998]);
csa_3018 csau_3018_i1266(tree_4[510041:507024],tree_4[513059:510042],tree_4[516077:513060],tree_5[341033:338016],tree_5[344051:341034]);
csa_3018 csau_3018_i1267(tree_4[519095:516078],tree_4[522113:519096],tree_4[525131:522114],tree_5[347069:344052],tree_5[350087:347070]);
csa_3018 csau_3018_i1268(tree_4[528149:525132],tree_4[531167:528150],tree_4[534185:531168],tree_5[353105:350088],tree_5[356123:353106]);
csa_3018 csau_3018_i1269(tree_4[537203:534186],tree_4[540221:537204],tree_4[543239:540222],tree_5[359141:356124],tree_5[362159:359142]);
csa_3018 csau_3018_i1270(tree_4[546257:543240],tree_4[549275:546258],tree_4[552293:549276],tree_5[365177:362160],tree_5[368195:365178]);
csa_3018 csau_3018_i1271(tree_4[555311:552294],tree_4[558329:555312],tree_4[561347:558330],tree_5[371213:368196],tree_5[374231:371214]);
csa_3018 csau_3018_i1272(tree_4[564365:561348],tree_4[567383:564366],tree_4[570401:567384],tree_5[377249:374232],tree_5[380267:377250]);
csa_3018 csau_3018_i1273(tree_4[573419:570402],tree_4[576437:573420],tree_4[579455:576438],tree_5[383285:380268],tree_5[386303:383286]);
csa_3018 csau_3018_i1274(tree_4[582473:579456],tree_4[585491:582474],tree_4[588509:585492],tree_5[389321:386304],tree_5[392339:389322]);
csa_3018 csau_3018_i1275(tree_4[591527:588510],tree_4[594545:591528],tree_4[597563:594546],tree_5[395357:392340],tree_5[398375:395358]);
csa_3018 csau_3018_i1276(tree_4[600581:597564],tree_4[603599:600582],tree_4[606617:603600],tree_5[401393:398376],tree_5[404411:401394]);
csa_3018 csau_3018_i1277(tree_4[609635:606618],tree_4[612653:609636],tree_4[615671:612654],tree_5[407429:404412],tree_5[410447:407430]);
csa_3018 csau_3018_i1278(tree_4[618689:615672],tree_4[621707:618690],tree_4[624725:621708],tree_5[413465:410448],tree_5[416483:413466]);
csa_3018 csau_3018_i1279(tree_4[627743:624726],tree_4[630761:627744],tree_4[633779:630762],tree_5[419501:416484],tree_5[422519:419502]);
csa_3018 csau_3018_i1280(tree_4[636797:633780],tree_4[639815:636798],tree_4[642833:639816],tree_5[425537:422520],tree_5[428555:425538]);
csa_3018 csau_3018_i1281(tree_4[645851:642834],tree_4[648869:645852],tree_4[651887:648870],tree_5[431573:428556],tree_5[434591:431574]);
csa_3018 csau_3018_i1282(tree_4[654905:651888],tree_4[657923:654906],tree_4[660941:657924],tree_5[437609:434592],tree_5[440627:437610]);
csa_3018 csau_3018_i1283(tree_4[663959:660942],tree_4[666977:663960],tree_4[669995:666978],tree_5[443645:440628],tree_5[446663:443646]);
csa_3018 csau_3018_i1284(tree_4[673013:669996],tree_4[676031:673014],tree_4[679049:676032],tree_5[449681:446664],tree_5[452699:449682]);
csa_3018 csau_3018_i1285(tree_4[682067:679050],tree_4[685085:682068],tree_4[688103:685086],tree_5[455717:452700],tree_5[458735:455718]);
csa_3018 csau_3018_i1286(tree_4[691121:688104],tree_4[694139:691122],tree_4[697157:694140],tree_5[461753:458736],tree_5[464771:461754]);
csa_3018 csau_3018_i1287(tree_4[700175:697158],tree_4[703193:700176],tree_4[706211:703194],tree_5[467789:464772],tree_5[470807:467790]);
csa_3018 csau_3018_i1288(tree_4[709229:706212],tree_4[712247:709230],tree_4[715265:712248],tree_5[473825:470808],tree_5[476843:473826]);
csa_3018 csau_3018_i1289(tree_4[718283:715266],tree_4[721301:718284],tree_4[724319:721302],tree_5[479861:476844],tree_5[482879:479862]);
csa_3018 csau_3018_i1290(tree_4[727337:724320],tree_4[730355:727338],tree_4[733373:730356],tree_5[485897:482880],tree_5[488915:485898]);
csa_3018 csau_3018_i1291(tree_4[736391:733374],tree_4[739409:736392],tree_4[742427:739410],tree_5[491933:488916],tree_5[494951:491934]);
csa_3018 csau_3018_i1292(tree_4[745445:742428],tree_4[748463:745446],tree_4[751481:748464],tree_5[497969:494952],tree_5[500987:497970]);
csa_3018 csau_3018_i1293(tree_4[754499:751482],tree_4[757517:754500],tree_4[760535:757518],tree_5[504005:500988],tree_5[507023:504006]);
csa_3018 csau_3018_i1294(tree_4[763553:760536],tree_4[766571:763554],tree_4[769589:766572],tree_5[510041:507024],tree_5[513059:510042]);
csa_3018 csau_3018_i1295(tree_4[772607:769590],tree_4[775625:772608],tree_4[778643:775626],tree_5[516077:513060],tree_5[519095:516078]);
csa_3018 csau_3018_i1296(tree_4[781661:778644],tree_4[784679:781662],tree_4[787697:784680],tree_5[522113:519096],tree_5[525131:522114]);
csa_3018 csau_3018_i1297(tree_4[790715:787698],tree_4[793733:790716],tree_4[796751:793734],tree_5[528149:525132],tree_5[531167:528150]);
csa_3018 csau_3018_i1298(tree_4[799769:796752],tree_4[802787:799770],tree_4[805805:802788],tree_5[534185:531168],tree_5[537203:534186]);
csa_3018 csau_3018_i1299(tree_4[808823:805806],tree_4[811841:808824],tree_4[814859:811842],tree_5[540221:537204],tree_5[543239:540222]);
csa_3018 csau_3018_i1300(tree_4[817877:814860],tree_4[820895:817878],tree_4[823913:820896],tree_5[546257:543240],tree_5[549275:546258]);
csa_3018 csau_3018_i1301(tree_4[826931:823914],tree_4[829949:826932],tree_4[832967:829950],tree_5[552293:549276],tree_5[555311:552294]);
csa_3018 csau_3018_i1302(tree_4[835985:832968],tree_4[839003:835986],tree_4[842021:839004],tree_5[558329:555312],tree_5[561347:558330]);
csa_3018 csau_3018_i1303(tree_4[845039:842022],tree_4[848057:845040],tree_4[851075:848058],tree_5[564365:561348],tree_5[567383:564366]);
csa_3018 csau_3018_i1304(tree_4[854093:851076],tree_4[857111:854094],tree_4[860129:857112],tree_5[570401:567384],tree_5[573419:570402]);
csa_3018 csau_3018_i1305(tree_4[863147:860130],tree_4[866165:863148],tree_4[869183:866166],tree_5[576437:573420],tree_5[579455:576438]);
csa_3018 csau_3018_i1306(tree_4[872201:869184],tree_4[875219:872202],tree_4[878237:875220],tree_5[582473:579456],tree_5[585491:582474]);
csa_3018 csau_3018_i1307(tree_4[881255:878238],tree_4[884273:881256],tree_4[887291:884274],tree_5[588509:585492],tree_5[591527:588510]);
csa_3018 csau_3018_i1308(tree_4[890309:887292],tree_4[893327:890310],tree_4[896345:893328],tree_5[594545:591528],tree_5[597563:594546]);
assign tree_5[600581:597564] = tree_4[899363:896346];
assign tree_5[603599:600582] = tree_4[902381:899364];
// layer-6
csa_3018 csau_3018_i1309(tree_5[3017:0],tree_5[6035:3018],tree_5[9053:6036],tree_6[3017:0],tree_6[6035:3018]);
csa_3018 csau_3018_i1310(tree_5[12071:9054],tree_5[15089:12072],tree_5[18107:15090],tree_6[9053:6036],tree_6[12071:9054]);
csa_3018 csau_3018_i1311(tree_5[21125:18108],tree_5[24143:21126],tree_5[27161:24144],tree_6[15089:12072],tree_6[18107:15090]);
csa_3018 csau_3018_i1312(tree_5[30179:27162],tree_5[33197:30180],tree_5[36215:33198],tree_6[21125:18108],tree_6[24143:21126]);
csa_3018 csau_3018_i1313(tree_5[39233:36216],tree_5[42251:39234],tree_5[45269:42252],tree_6[27161:24144],tree_6[30179:27162]);
csa_3018 csau_3018_i1314(tree_5[48287:45270],tree_5[51305:48288],tree_5[54323:51306],tree_6[33197:30180],tree_6[36215:33198]);
csa_3018 csau_3018_i1315(tree_5[57341:54324],tree_5[60359:57342],tree_5[63377:60360],tree_6[39233:36216],tree_6[42251:39234]);
csa_3018 csau_3018_i1316(tree_5[66395:63378],tree_5[69413:66396],tree_5[72431:69414],tree_6[45269:42252],tree_6[48287:45270]);
csa_3018 csau_3018_i1317(tree_5[75449:72432],tree_5[78467:75450],tree_5[81485:78468],tree_6[51305:48288],tree_6[54323:51306]);
csa_3018 csau_3018_i1318(tree_5[84503:81486],tree_5[87521:84504],tree_5[90539:87522],tree_6[57341:54324],tree_6[60359:57342]);
csa_3018 csau_3018_i1319(tree_5[93557:90540],tree_5[96575:93558],tree_5[99593:96576],tree_6[63377:60360],tree_6[66395:63378]);
csa_3018 csau_3018_i1320(tree_5[102611:99594],tree_5[105629:102612],tree_5[108647:105630],tree_6[69413:66396],tree_6[72431:69414]);
csa_3018 csau_3018_i1321(tree_5[111665:108648],tree_5[114683:111666],tree_5[117701:114684],tree_6[75449:72432],tree_6[78467:75450]);
csa_3018 csau_3018_i1322(tree_5[120719:117702],tree_5[123737:120720],tree_5[126755:123738],tree_6[81485:78468],tree_6[84503:81486]);
csa_3018 csau_3018_i1323(tree_5[129773:126756],tree_5[132791:129774],tree_5[135809:132792],tree_6[87521:84504],tree_6[90539:87522]);
csa_3018 csau_3018_i1324(tree_5[138827:135810],tree_5[141845:138828],tree_5[144863:141846],tree_6[93557:90540],tree_6[96575:93558]);
csa_3018 csau_3018_i1325(tree_5[147881:144864],tree_5[150899:147882],tree_5[153917:150900],tree_6[99593:96576],tree_6[102611:99594]);
csa_3018 csau_3018_i1326(tree_5[156935:153918],tree_5[159953:156936],tree_5[162971:159954],tree_6[105629:102612],tree_6[108647:105630]);
csa_3018 csau_3018_i1327(tree_5[165989:162972],tree_5[169007:165990],tree_5[172025:169008],tree_6[111665:108648],tree_6[114683:111666]);
csa_3018 csau_3018_i1328(tree_5[175043:172026],tree_5[178061:175044],tree_5[181079:178062],tree_6[117701:114684],tree_6[120719:117702]);
csa_3018 csau_3018_i1329(tree_5[184097:181080],tree_5[187115:184098],tree_5[190133:187116],tree_6[123737:120720],tree_6[126755:123738]);
csa_3018 csau_3018_i1330(tree_5[193151:190134],tree_5[196169:193152],tree_5[199187:196170],tree_6[129773:126756],tree_6[132791:129774]);
csa_3018 csau_3018_i1331(tree_5[202205:199188],tree_5[205223:202206],tree_5[208241:205224],tree_6[135809:132792],tree_6[138827:135810]);
csa_3018 csau_3018_i1332(tree_5[211259:208242],tree_5[214277:211260],tree_5[217295:214278],tree_6[141845:138828],tree_6[144863:141846]);
csa_3018 csau_3018_i1333(tree_5[220313:217296],tree_5[223331:220314],tree_5[226349:223332],tree_6[147881:144864],tree_6[150899:147882]);
csa_3018 csau_3018_i1334(tree_5[229367:226350],tree_5[232385:229368],tree_5[235403:232386],tree_6[153917:150900],tree_6[156935:153918]);
csa_3018 csau_3018_i1335(tree_5[238421:235404],tree_5[241439:238422],tree_5[244457:241440],tree_6[159953:156936],tree_6[162971:159954]);
csa_3018 csau_3018_i1336(tree_5[247475:244458],tree_5[250493:247476],tree_5[253511:250494],tree_6[165989:162972],tree_6[169007:165990]);
csa_3018 csau_3018_i1337(tree_5[256529:253512],tree_5[259547:256530],tree_5[262565:259548],tree_6[172025:169008],tree_6[175043:172026]);
csa_3018 csau_3018_i1338(tree_5[265583:262566],tree_5[268601:265584],tree_5[271619:268602],tree_6[178061:175044],tree_6[181079:178062]);
csa_3018 csau_3018_i1339(tree_5[274637:271620],tree_5[277655:274638],tree_5[280673:277656],tree_6[184097:181080],tree_6[187115:184098]);
csa_3018 csau_3018_i1340(tree_5[283691:280674],tree_5[286709:283692],tree_5[289727:286710],tree_6[190133:187116],tree_6[193151:190134]);
csa_3018 csau_3018_i1341(tree_5[292745:289728],tree_5[295763:292746],tree_5[298781:295764],tree_6[196169:193152],tree_6[199187:196170]);
csa_3018 csau_3018_i1342(tree_5[301799:298782],tree_5[304817:301800],tree_5[307835:304818],tree_6[202205:199188],tree_6[205223:202206]);
csa_3018 csau_3018_i1343(tree_5[310853:307836],tree_5[313871:310854],tree_5[316889:313872],tree_6[208241:205224],tree_6[211259:208242]);
csa_3018 csau_3018_i1344(tree_5[319907:316890],tree_5[322925:319908],tree_5[325943:322926],tree_6[214277:211260],tree_6[217295:214278]);
csa_3018 csau_3018_i1345(tree_5[328961:325944],tree_5[331979:328962],tree_5[334997:331980],tree_6[220313:217296],tree_6[223331:220314]);
csa_3018 csau_3018_i1346(tree_5[338015:334998],tree_5[341033:338016],tree_5[344051:341034],tree_6[226349:223332],tree_6[229367:226350]);
csa_3018 csau_3018_i1347(tree_5[347069:344052],tree_5[350087:347070],tree_5[353105:350088],tree_6[232385:229368],tree_6[235403:232386]);
csa_3018 csau_3018_i1348(tree_5[356123:353106],tree_5[359141:356124],tree_5[362159:359142],tree_6[238421:235404],tree_6[241439:238422]);
csa_3018 csau_3018_i1349(tree_5[365177:362160],tree_5[368195:365178],tree_5[371213:368196],tree_6[244457:241440],tree_6[247475:244458]);
csa_3018 csau_3018_i1350(tree_5[374231:371214],tree_5[377249:374232],tree_5[380267:377250],tree_6[250493:247476],tree_6[253511:250494]);
csa_3018 csau_3018_i1351(tree_5[383285:380268],tree_5[386303:383286],tree_5[389321:386304],tree_6[256529:253512],tree_6[259547:256530]);
csa_3018 csau_3018_i1352(tree_5[392339:389322],tree_5[395357:392340],tree_5[398375:395358],tree_6[262565:259548],tree_6[265583:262566]);
csa_3018 csau_3018_i1353(tree_5[401393:398376],tree_5[404411:401394],tree_5[407429:404412],tree_6[268601:265584],tree_6[271619:268602]);
csa_3018 csau_3018_i1354(tree_5[410447:407430],tree_5[413465:410448],tree_5[416483:413466],tree_6[274637:271620],tree_6[277655:274638]);
csa_3018 csau_3018_i1355(tree_5[419501:416484],tree_5[422519:419502],tree_5[425537:422520],tree_6[280673:277656],tree_6[283691:280674]);
csa_3018 csau_3018_i1356(tree_5[428555:425538],tree_5[431573:428556],tree_5[434591:431574],tree_6[286709:283692],tree_6[289727:286710]);
csa_3018 csau_3018_i1357(tree_5[437609:434592],tree_5[440627:437610],tree_5[443645:440628],tree_6[292745:289728],tree_6[295763:292746]);
csa_3018 csau_3018_i1358(tree_5[446663:443646],tree_5[449681:446664],tree_5[452699:449682],tree_6[298781:295764],tree_6[301799:298782]);
csa_3018 csau_3018_i1359(tree_5[455717:452700],tree_5[458735:455718],tree_5[461753:458736],tree_6[304817:301800],tree_6[307835:304818]);
csa_3018 csau_3018_i1360(tree_5[464771:461754],tree_5[467789:464772],tree_5[470807:467790],tree_6[310853:307836],tree_6[313871:310854]);
csa_3018 csau_3018_i1361(tree_5[473825:470808],tree_5[476843:473826],tree_5[479861:476844],tree_6[316889:313872],tree_6[319907:316890]);
csa_3018 csau_3018_i1362(tree_5[482879:479862],tree_5[485897:482880],tree_5[488915:485898],tree_6[322925:319908],tree_6[325943:322926]);
csa_3018 csau_3018_i1363(tree_5[491933:488916],tree_5[494951:491934],tree_5[497969:494952],tree_6[328961:325944],tree_6[331979:328962]);
csa_3018 csau_3018_i1364(tree_5[500987:497970],tree_5[504005:500988],tree_5[507023:504006],tree_6[334997:331980],tree_6[338015:334998]);
csa_3018 csau_3018_i1365(tree_5[510041:507024],tree_5[513059:510042],tree_5[516077:513060],tree_6[341033:338016],tree_6[344051:341034]);
csa_3018 csau_3018_i1366(tree_5[519095:516078],tree_5[522113:519096],tree_5[525131:522114],tree_6[347069:344052],tree_6[350087:347070]);
csa_3018 csau_3018_i1367(tree_5[528149:525132],tree_5[531167:528150],tree_5[534185:531168],tree_6[353105:350088],tree_6[356123:353106]);
csa_3018 csau_3018_i1368(tree_5[537203:534186],tree_5[540221:537204],tree_5[543239:540222],tree_6[359141:356124],tree_6[362159:359142]);
csa_3018 csau_3018_i1369(tree_5[546257:543240],tree_5[549275:546258],tree_5[552293:549276],tree_6[365177:362160],tree_6[368195:365178]);
csa_3018 csau_3018_i1370(tree_5[555311:552294],tree_5[558329:555312],tree_5[561347:558330],tree_6[371213:368196],tree_6[374231:371214]);
csa_3018 csau_3018_i1371(tree_5[564365:561348],tree_5[567383:564366],tree_5[570401:567384],tree_6[377249:374232],tree_6[380267:377250]);
csa_3018 csau_3018_i1372(tree_5[573419:570402],tree_5[576437:573420],tree_5[579455:576438],tree_6[383285:380268],tree_6[386303:383286]);
csa_3018 csau_3018_i1373(tree_5[582473:579456],tree_5[585491:582474],tree_5[588509:585492],tree_6[389321:386304],tree_6[392339:389322]);
csa_3018 csau_3018_i1374(tree_5[591527:588510],tree_5[594545:591528],tree_5[597563:594546],tree_6[395357:392340],tree_6[398375:395358]);
assign tree_6[401393:398376] = tree_5[600581:597564];
assign tree_6[404411:401394] = tree_5[603599:600582];
// layer-7
csa_3018 csau_3018_i1375(tree_6[3017:0],tree_6[6035:3018],tree_6[9053:6036],tree_7[3017:0],tree_7[6035:3018]);
csa_3018 csau_3018_i1376(tree_6[12071:9054],tree_6[15089:12072],tree_6[18107:15090],tree_7[9053:6036],tree_7[12071:9054]);
csa_3018 csau_3018_i1377(tree_6[21125:18108],tree_6[24143:21126],tree_6[27161:24144],tree_7[15089:12072],tree_7[18107:15090]);
csa_3018 csau_3018_i1378(tree_6[30179:27162],tree_6[33197:30180],tree_6[36215:33198],tree_7[21125:18108],tree_7[24143:21126]);
csa_3018 csau_3018_i1379(tree_6[39233:36216],tree_6[42251:39234],tree_6[45269:42252],tree_7[27161:24144],tree_7[30179:27162]);
csa_3018 csau_3018_i1380(tree_6[48287:45270],tree_6[51305:48288],tree_6[54323:51306],tree_7[33197:30180],tree_7[36215:33198]);
csa_3018 csau_3018_i1381(tree_6[57341:54324],tree_6[60359:57342],tree_6[63377:60360],tree_7[39233:36216],tree_7[42251:39234]);
csa_3018 csau_3018_i1382(tree_6[66395:63378],tree_6[69413:66396],tree_6[72431:69414],tree_7[45269:42252],tree_7[48287:45270]);
csa_3018 csau_3018_i1383(tree_6[75449:72432],tree_6[78467:75450],tree_6[81485:78468],tree_7[51305:48288],tree_7[54323:51306]);
csa_3018 csau_3018_i1384(tree_6[84503:81486],tree_6[87521:84504],tree_6[90539:87522],tree_7[57341:54324],tree_7[60359:57342]);
csa_3018 csau_3018_i1385(tree_6[93557:90540],tree_6[96575:93558],tree_6[99593:96576],tree_7[63377:60360],tree_7[66395:63378]);
csa_3018 csau_3018_i1386(tree_6[102611:99594],tree_6[105629:102612],tree_6[108647:105630],tree_7[69413:66396],tree_7[72431:69414]);
csa_3018 csau_3018_i1387(tree_6[111665:108648],tree_6[114683:111666],tree_6[117701:114684],tree_7[75449:72432],tree_7[78467:75450]);
csa_3018 csau_3018_i1388(tree_6[120719:117702],tree_6[123737:120720],tree_6[126755:123738],tree_7[81485:78468],tree_7[84503:81486]);
csa_3018 csau_3018_i1389(tree_6[129773:126756],tree_6[132791:129774],tree_6[135809:132792],tree_7[87521:84504],tree_7[90539:87522]);
csa_3018 csau_3018_i1390(tree_6[138827:135810],tree_6[141845:138828],tree_6[144863:141846],tree_7[93557:90540],tree_7[96575:93558]);
csa_3018 csau_3018_i1391(tree_6[147881:144864],tree_6[150899:147882],tree_6[153917:150900],tree_7[99593:96576],tree_7[102611:99594]);
csa_3018 csau_3018_i1392(tree_6[156935:153918],tree_6[159953:156936],tree_6[162971:159954],tree_7[105629:102612],tree_7[108647:105630]);
csa_3018 csau_3018_i1393(tree_6[165989:162972],tree_6[169007:165990],tree_6[172025:169008],tree_7[111665:108648],tree_7[114683:111666]);
csa_3018 csau_3018_i1394(tree_6[175043:172026],tree_6[178061:175044],tree_6[181079:178062],tree_7[117701:114684],tree_7[120719:117702]);
csa_3018 csau_3018_i1395(tree_6[184097:181080],tree_6[187115:184098],tree_6[190133:187116],tree_7[123737:120720],tree_7[126755:123738]);
csa_3018 csau_3018_i1396(tree_6[193151:190134],tree_6[196169:193152],tree_6[199187:196170],tree_7[129773:126756],tree_7[132791:129774]);
csa_3018 csau_3018_i1397(tree_6[202205:199188],tree_6[205223:202206],tree_6[208241:205224],tree_7[135809:132792],tree_7[138827:135810]);
csa_3018 csau_3018_i1398(tree_6[211259:208242],tree_6[214277:211260],tree_6[217295:214278],tree_7[141845:138828],tree_7[144863:141846]);
csa_3018 csau_3018_i1399(tree_6[220313:217296],tree_6[223331:220314],tree_6[226349:223332],tree_7[147881:144864],tree_7[150899:147882]);
csa_3018 csau_3018_i1400(tree_6[229367:226350],tree_6[232385:229368],tree_6[235403:232386],tree_7[153917:150900],tree_7[156935:153918]);
csa_3018 csau_3018_i1401(tree_6[238421:235404],tree_6[241439:238422],tree_6[244457:241440],tree_7[159953:156936],tree_7[162971:159954]);
csa_3018 csau_3018_i1402(tree_6[247475:244458],tree_6[250493:247476],tree_6[253511:250494],tree_7[165989:162972],tree_7[169007:165990]);
csa_3018 csau_3018_i1403(tree_6[256529:253512],tree_6[259547:256530],tree_6[262565:259548],tree_7[172025:169008],tree_7[175043:172026]);
csa_3018 csau_3018_i1404(tree_6[265583:262566],tree_6[268601:265584],tree_6[271619:268602],tree_7[178061:175044],tree_7[181079:178062]);
csa_3018 csau_3018_i1405(tree_6[274637:271620],tree_6[277655:274638],tree_6[280673:277656],tree_7[184097:181080],tree_7[187115:184098]);
csa_3018 csau_3018_i1406(tree_6[283691:280674],tree_6[286709:283692],tree_6[289727:286710],tree_7[190133:187116],tree_7[193151:190134]);
csa_3018 csau_3018_i1407(tree_6[292745:289728],tree_6[295763:292746],tree_6[298781:295764],tree_7[196169:193152],tree_7[199187:196170]);
csa_3018 csau_3018_i1408(tree_6[301799:298782],tree_6[304817:301800],tree_6[307835:304818],tree_7[202205:199188],tree_7[205223:202206]);
csa_3018 csau_3018_i1409(tree_6[310853:307836],tree_6[313871:310854],tree_6[316889:313872],tree_7[208241:205224],tree_7[211259:208242]);
csa_3018 csau_3018_i1410(tree_6[319907:316890],tree_6[322925:319908],tree_6[325943:322926],tree_7[214277:211260],tree_7[217295:214278]);
csa_3018 csau_3018_i1411(tree_6[328961:325944],tree_6[331979:328962],tree_6[334997:331980],tree_7[220313:217296],tree_7[223331:220314]);
csa_3018 csau_3018_i1412(tree_6[338015:334998],tree_6[341033:338016],tree_6[344051:341034],tree_7[226349:223332],tree_7[229367:226350]);
csa_3018 csau_3018_i1413(tree_6[347069:344052],tree_6[350087:347070],tree_6[353105:350088],tree_7[232385:229368],tree_7[235403:232386]);
csa_3018 csau_3018_i1414(tree_6[356123:353106],tree_6[359141:356124],tree_6[362159:359142],tree_7[238421:235404],tree_7[241439:238422]);
csa_3018 csau_3018_i1415(tree_6[365177:362160],tree_6[368195:365178],tree_6[371213:368196],tree_7[244457:241440],tree_7[247475:244458]);
csa_3018 csau_3018_i1416(tree_6[374231:371214],tree_6[377249:374232],tree_6[380267:377250],tree_7[250493:247476],tree_7[253511:250494]);
csa_3018 csau_3018_i1417(tree_6[383285:380268],tree_6[386303:383286],tree_6[389321:386304],tree_7[256529:253512],tree_7[259547:256530]);
csa_3018 csau_3018_i1418(tree_6[392339:389322],tree_6[395357:392340],tree_6[398375:395358],tree_7[262565:259548],tree_7[265583:262566]);
assign tree_7[268601:265584] = tree_6[401393:398376];
assign tree_7[271619:268602] = tree_6[404411:401394];
// layer-8
csa_3018 csau_3018_i1419(tree_7[3017:0],tree_7[6035:3018],tree_7[9053:6036],tree_8[3017:0],tree_8[6035:3018]);
csa_3018 csau_3018_i1420(tree_7[12071:9054],tree_7[15089:12072],tree_7[18107:15090],tree_8[9053:6036],tree_8[12071:9054]);
csa_3018 csau_3018_i1421(tree_7[21125:18108],tree_7[24143:21126],tree_7[27161:24144],tree_8[15089:12072],tree_8[18107:15090]);
csa_3018 csau_3018_i1422(tree_7[30179:27162],tree_7[33197:30180],tree_7[36215:33198],tree_8[21125:18108],tree_8[24143:21126]);
csa_3018 csau_3018_i1423(tree_7[39233:36216],tree_7[42251:39234],tree_7[45269:42252],tree_8[27161:24144],tree_8[30179:27162]);
csa_3018 csau_3018_i1424(tree_7[48287:45270],tree_7[51305:48288],tree_7[54323:51306],tree_8[33197:30180],tree_8[36215:33198]);
csa_3018 csau_3018_i1425(tree_7[57341:54324],tree_7[60359:57342],tree_7[63377:60360],tree_8[39233:36216],tree_8[42251:39234]);
csa_3018 csau_3018_i1426(tree_7[66395:63378],tree_7[69413:66396],tree_7[72431:69414],tree_8[45269:42252],tree_8[48287:45270]);
csa_3018 csau_3018_i1427(tree_7[75449:72432],tree_7[78467:75450],tree_7[81485:78468],tree_8[51305:48288],tree_8[54323:51306]);
csa_3018 csau_3018_i1428(tree_7[84503:81486],tree_7[87521:84504],tree_7[90539:87522],tree_8[57341:54324],tree_8[60359:57342]);
csa_3018 csau_3018_i1429(tree_7[93557:90540],tree_7[96575:93558],tree_7[99593:96576],tree_8[63377:60360],tree_8[66395:63378]);
csa_3018 csau_3018_i1430(tree_7[102611:99594],tree_7[105629:102612],tree_7[108647:105630],tree_8[69413:66396],tree_8[72431:69414]);
csa_3018 csau_3018_i1431(tree_7[111665:108648],tree_7[114683:111666],tree_7[117701:114684],tree_8[75449:72432],tree_8[78467:75450]);
csa_3018 csau_3018_i1432(tree_7[120719:117702],tree_7[123737:120720],tree_7[126755:123738],tree_8[81485:78468],tree_8[84503:81486]);
csa_3018 csau_3018_i1433(tree_7[129773:126756],tree_7[132791:129774],tree_7[135809:132792],tree_8[87521:84504],tree_8[90539:87522]);
csa_3018 csau_3018_i1434(tree_7[138827:135810],tree_7[141845:138828],tree_7[144863:141846],tree_8[93557:90540],tree_8[96575:93558]);
csa_3018 csau_3018_i1435(tree_7[147881:144864],tree_7[150899:147882],tree_7[153917:150900],tree_8[99593:96576],tree_8[102611:99594]);
csa_3018 csau_3018_i1436(tree_7[156935:153918],tree_7[159953:156936],tree_7[162971:159954],tree_8[105629:102612],tree_8[108647:105630]);
csa_3018 csau_3018_i1437(tree_7[165989:162972],tree_7[169007:165990],tree_7[172025:169008],tree_8[111665:108648],tree_8[114683:111666]);
csa_3018 csau_3018_i1438(tree_7[175043:172026],tree_7[178061:175044],tree_7[181079:178062],tree_8[117701:114684],tree_8[120719:117702]);
csa_3018 csau_3018_i1439(tree_7[184097:181080],tree_7[187115:184098],tree_7[190133:187116],tree_8[123737:120720],tree_8[126755:123738]);
csa_3018 csau_3018_i1440(tree_7[193151:190134],tree_7[196169:193152],tree_7[199187:196170],tree_8[129773:126756],tree_8[132791:129774]);
csa_3018 csau_3018_i1441(tree_7[202205:199188],tree_7[205223:202206],tree_7[208241:205224],tree_8[135809:132792],tree_8[138827:135810]);
csa_3018 csau_3018_i1442(tree_7[211259:208242],tree_7[214277:211260],tree_7[217295:214278],tree_8[141845:138828],tree_8[144863:141846]);
csa_3018 csau_3018_i1443(tree_7[220313:217296],tree_7[223331:220314],tree_7[226349:223332],tree_8[147881:144864],tree_8[150899:147882]);
csa_3018 csau_3018_i1444(tree_7[229367:226350],tree_7[232385:229368],tree_7[235403:232386],tree_8[153917:150900],tree_8[156935:153918]);
csa_3018 csau_3018_i1445(tree_7[238421:235404],tree_7[241439:238422],tree_7[244457:241440],tree_8[159953:156936],tree_8[162971:159954]);
csa_3018 csau_3018_i1446(tree_7[247475:244458],tree_7[250493:247476],tree_7[253511:250494],tree_8[165989:162972],tree_8[169007:165990]);
csa_3018 csau_3018_i1447(tree_7[256529:253512],tree_7[259547:256530],tree_7[262565:259548],tree_8[172025:169008],tree_8[175043:172026]);
csa_3018 csau_3018_i1448(tree_7[265583:262566],tree_7[268601:265584],tree_7[271619:268602],tree_8[178061:175044],tree_8[181079:178062]);
// layer-9
csa_3018 csau_3018_i1449(tree_8[3017:0],tree_8[6035:3018],tree_8[9053:6036],tree_9[3017:0],tree_9[6035:3018]);
csa_3018 csau_3018_i1450(tree_8[12071:9054],tree_8[15089:12072],tree_8[18107:15090],tree_9[9053:6036],tree_9[12071:9054]);
csa_3018 csau_3018_i1451(tree_8[21125:18108],tree_8[24143:21126],tree_8[27161:24144],tree_9[15089:12072],tree_9[18107:15090]);
csa_3018 csau_3018_i1452(tree_8[30179:27162],tree_8[33197:30180],tree_8[36215:33198],tree_9[21125:18108],tree_9[24143:21126]);
csa_3018 csau_3018_i1453(tree_8[39233:36216],tree_8[42251:39234],tree_8[45269:42252],tree_9[27161:24144],tree_9[30179:27162]);
csa_3018 csau_3018_i1454(tree_8[48287:45270],tree_8[51305:48288],tree_8[54323:51306],tree_9[33197:30180],tree_9[36215:33198]);
csa_3018 csau_3018_i1455(tree_8[57341:54324],tree_8[60359:57342],tree_8[63377:60360],tree_9[39233:36216],tree_9[42251:39234]);
csa_3018 csau_3018_i1456(tree_8[66395:63378],tree_8[69413:66396],tree_8[72431:69414],tree_9[45269:42252],tree_9[48287:45270]);
csa_3018 csau_3018_i1457(tree_8[75449:72432],tree_8[78467:75450],tree_8[81485:78468],tree_9[51305:48288],tree_9[54323:51306]);
csa_3018 csau_3018_i1458(tree_8[84503:81486],tree_8[87521:84504],tree_8[90539:87522],tree_9[57341:54324],tree_9[60359:57342]);
csa_3018 csau_3018_i1459(tree_8[93557:90540],tree_8[96575:93558],tree_8[99593:96576],tree_9[63377:60360],tree_9[66395:63378]);
csa_3018 csau_3018_i1460(tree_8[102611:99594],tree_8[105629:102612],tree_8[108647:105630],tree_9[69413:66396],tree_9[72431:69414]);
csa_3018 csau_3018_i1461(tree_8[111665:108648],tree_8[114683:111666],tree_8[117701:114684],tree_9[75449:72432],tree_9[78467:75450]);
csa_3018 csau_3018_i1462(tree_8[120719:117702],tree_8[123737:120720],tree_8[126755:123738],tree_9[81485:78468],tree_9[84503:81486]);
csa_3018 csau_3018_i1463(tree_8[129773:126756],tree_8[132791:129774],tree_8[135809:132792],tree_9[87521:84504],tree_9[90539:87522]);
csa_3018 csau_3018_i1464(tree_8[138827:135810],tree_8[141845:138828],tree_8[144863:141846],tree_9[93557:90540],tree_9[96575:93558]);
csa_3018 csau_3018_i1465(tree_8[147881:144864],tree_8[150899:147882],tree_8[153917:150900],tree_9[99593:96576],tree_9[102611:99594]);
csa_3018 csau_3018_i1466(tree_8[156935:153918],tree_8[159953:156936],tree_8[162971:159954],tree_9[105629:102612],tree_9[108647:105630]);
csa_3018 csau_3018_i1467(tree_8[165989:162972],tree_8[169007:165990],tree_8[172025:169008],tree_9[111665:108648],tree_9[114683:111666]);
csa_3018 csau_3018_i1468(tree_8[175043:172026],tree_8[178061:175044],tree_8[181079:178062],tree_9[117701:114684],tree_9[120719:117702]);
// layer-10
csa_3018 csau_3018_i1469(tree_9[3017:0],tree_9[6035:3018],tree_9[9053:6036],tree_10[3017:0],tree_10[6035:3018]);
csa_3018 csau_3018_i1470(tree_9[12071:9054],tree_9[15089:12072],tree_9[18107:15090],tree_10[9053:6036],tree_10[12071:9054]);
csa_3018 csau_3018_i1471(tree_9[21125:18108],tree_9[24143:21126],tree_9[27161:24144],tree_10[15089:12072],tree_10[18107:15090]);
csa_3018 csau_3018_i1472(tree_9[30179:27162],tree_9[33197:30180],tree_9[36215:33198],tree_10[21125:18108],tree_10[24143:21126]);
csa_3018 csau_3018_i1473(tree_9[39233:36216],tree_9[42251:39234],tree_9[45269:42252],tree_10[27161:24144],tree_10[30179:27162]);
csa_3018 csau_3018_i1474(tree_9[48287:45270],tree_9[51305:48288],tree_9[54323:51306],tree_10[33197:30180],tree_10[36215:33198]);
csa_3018 csau_3018_i1475(tree_9[57341:54324],tree_9[60359:57342],tree_9[63377:60360],tree_10[39233:36216],tree_10[42251:39234]);
csa_3018 csau_3018_i1476(tree_9[66395:63378],tree_9[69413:66396],tree_9[72431:69414],tree_10[45269:42252],tree_10[48287:45270]);
csa_3018 csau_3018_i1477(tree_9[75449:72432],tree_9[78467:75450],tree_9[81485:78468],tree_10[51305:48288],tree_10[54323:51306]);
csa_3018 csau_3018_i1478(tree_9[84503:81486],tree_9[87521:84504],tree_9[90539:87522],tree_10[57341:54324],tree_10[60359:57342]);
csa_3018 csau_3018_i1479(tree_9[93557:90540],tree_9[96575:93558],tree_9[99593:96576],tree_10[63377:60360],tree_10[66395:63378]);
csa_3018 csau_3018_i1480(tree_9[102611:99594],tree_9[105629:102612],tree_9[108647:105630],tree_10[69413:66396],tree_10[72431:69414]);
csa_3018 csau_3018_i1481(tree_9[111665:108648],tree_9[114683:111666],tree_9[117701:114684],tree_10[75449:72432],tree_10[78467:75450]);
assign tree_10[81485:78468] = tree_9[120719:117702];
// layer-11
csa_3018 csau_3018_i1482(tree_10[3017:0],tree_10[6035:3018],tree_10[9053:6036],tree_11[3017:0],tree_11[6035:3018]);
csa_3018 csau_3018_i1483(tree_10[12071:9054],tree_10[15089:12072],tree_10[18107:15090],tree_11[9053:6036],tree_11[12071:9054]);
csa_3018 csau_3018_i1484(tree_10[21125:18108],tree_10[24143:21126],tree_10[27161:24144],tree_11[15089:12072],tree_11[18107:15090]);
csa_3018 csau_3018_i1485(tree_10[30179:27162],tree_10[33197:30180],tree_10[36215:33198],tree_11[21125:18108],tree_11[24143:21126]);
csa_3018 csau_3018_i1486(tree_10[39233:36216],tree_10[42251:39234],tree_10[45269:42252],tree_11[27161:24144],tree_11[30179:27162]);
csa_3018 csau_3018_i1487(tree_10[48287:45270],tree_10[51305:48288],tree_10[54323:51306],tree_11[33197:30180],tree_11[36215:33198]);
csa_3018 csau_3018_i1488(tree_10[57341:54324],tree_10[60359:57342],tree_10[63377:60360],tree_11[39233:36216],tree_11[42251:39234]);
csa_3018 csau_3018_i1489(tree_10[66395:63378],tree_10[69413:66396],tree_10[72431:69414],tree_11[45269:42252],tree_11[48287:45270]);
csa_3018 csau_3018_i1490(tree_10[75449:72432],tree_10[78467:75450],tree_10[81485:78468],tree_11[51305:48288],tree_11[54323:51306]);
// layer-12
csa_3018 csau_3018_i1491(tree_11[3017:0],tree_11[6035:3018],tree_11[9053:6036],tree_12[3017:0],tree_12[6035:3018]);
csa_3018 csau_3018_i1492(tree_11[12071:9054],tree_11[15089:12072],tree_11[18107:15090],tree_12[9053:6036],tree_12[12071:9054]);
csa_3018 csau_3018_i1493(tree_11[21125:18108],tree_11[24143:21126],tree_11[27161:24144],tree_12[15089:12072],tree_12[18107:15090]);
csa_3018 csau_3018_i1494(tree_11[30179:27162],tree_11[33197:30180],tree_11[36215:33198],tree_12[21125:18108],tree_12[24143:21126]);
csa_3018 csau_3018_i1495(tree_11[39233:36216],tree_11[42251:39234],tree_11[45269:42252],tree_12[27161:24144],tree_12[30179:27162]);
csa_3018 csau_3018_i1496(tree_11[48287:45270],tree_11[51305:48288],tree_11[54323:51306],tree_12[33197:30180],tree_12[36215:33198]);
// layer-13
csa_3018 csau_3018_i1497(tree_12[3017:0],tree_12[6035:3018],tree_12[9053:6036],tree_13[3017:0],tree_13[6035:3018]);
csa_3018 csau_3018_i1498(tree_12[12071:9054],tree_12[15089:12072],tree_12[18107:15090],tree_13[9053:6036],tree_13[12071:9054]);
csa_3018 csau_3018_i1499(tree_12[21125:18108],tree_12[24143:21126],tree_12[27161:24144],tree_13[15089:12072],tree_13[18107:15090]);
csa_3018 csau_3018_i1500(tree_12[30179:27162],tree_12[33197:30180],tree_12[36215:33198],tree_13[21125:18108],tree_13[24143:21126]);
// layer-14
csa_3018 csau_3018_i1501(tree_13[3017:0],tree_13[6035:3018],tree_13[9053:6036],tree_14[3017:0],tree_14[6035:3018]);
csa_3018 csau_3018_i1502(tree_13[12071:9054],tree_13[15089:12072],tree_13[18107:15090],tree_14[9053:6036],tree_14[12071:9054]);
assign tree_14[15089:12072] = tree_13[21125:18108];
assign tree_14[18107:15090] = tree_13[24143:21126];
// layer-15
csa_3018 csau_3018_i1503(tree_14[3017:0],tree_14[6035:3018],tree_14[9053:6036],tree_15[3017:0],tree_15[6035:3018]);
csa_3018 csau_3018_i1504(tree_14[12071:9054],tree_14[15089:12072],tree_14[18107:15090],tree_15[9053:6036],tree_15[12071:9054]);
// layer-16
csa_3018 csau_3018_i1505(tree_15[3017:0],tree_15[6035:3018],tree_15[9053:6036],tree_16[3017:0],tree_16[6035:3018]);
assign tree_16[9053:6036] = tree_15[12071:9054];
// layer-17
csa_3018 csau_3018_i1506(tree_16[3017:0],tree_16[6035:3018],tree_16[9053:6036],tree_17[3017:0],tree_17[6035:3018]);

// final assignment
assign B_0 = tree_17[3017:0];
assign B_1 = tree_17[6035:3018];

endmodule
