
module red_part1_43x43(
    input [81:0] a_c,a_s,
    input [42:0] p_prime,
    output [1848:0] b_c,b_s // lines are appended together
);
    
wire [42:0] c_w_0, s_w_0;
wire [42:0] c_w_1, s_w_1;
wire [42:0] c_w_2, s_w_2;
wire [42:0] c_w_3, s_w_3;
wire [42:0] c_w_4, s_w_4;
wire [42:0] c_w_5, s_w_5;
wire [42:0] c_w_6, s_w_6;
wire [42:0] c_w_7, s_w_7;
wire [42:0] c_w_8, s_w_8;
wire [42:0] c_w_9, s_w_9;
wire [42:0] c_w_10, s_w_10;
wire [42:0] c_w_11, s_w_11;
wire [42:0] c_w_12, s_w_12;
wire [42:0] c_w_13, s_w_13;
wire [42:0] c_w_14, s_w_14;
wire [42:0] c_w_15, s_w_15;
wire [42:0] c_w_16, s_w_16;
wire [42:0] c_w_17, s_w_17;
wire [42:0] c_w_18, s_w_18;
wire [42:0] c_w_19, s_w_19;
wire [42:0] c_w_20, s_w_20;
wire [42:0] c_w_21, s_w_21;
wire [42:0] c_w_22, s_w_22;
wire [42:0] c_w_23, s_w_23;
wire [42:0] c_w_24, s_w_24;
wire [42:0] c_w_25, s_w_25;
wire [42:0] c_w_26, s_w_26;
wire [42:0] c_w_27, s_w_27;
wire [42:0] c_w_28, s_w_28;
wire [42:0] c_w_29, s_w_29;
wire [42:0] c_w_30, s_w_30;
wire [42:0] c_w_31, s_w_31;
wire [42:0] c_w_32, s_w_32;
wire [42:0] c_w_33, s_w_33;
wire [42:0] c_w_34, s_w_34;
wire [42:0] c_w_35, s_w_35;
wire [42:0] c_w_36, s_w_36;
wire [42:0] c_w_37, s_w_37;
wire [42:0] c_w_38, s_w_38;
wire [42:0] c_w_39, s_w_39;
wire [42:0] c_w_40, s_w_40;
wire [42:0] c_w_41, s_w_41;
wire [42:0] c_w_42, s_w_42;
    
AND_array_43 AND_array_43_c0({a_c[42:0]},p_prime[0],c_w_0);
AND_array_43 AND_array_43_s0({a_s[42:0]},p_prime[0],s_w_0);
AND_array_43 AND_array_43_c1({a_c[41:0],1'd0},p_prime[1],c_w_1);
AND_array_43 AND_array_43_s1({a_s[41:0],1'd0},p_prime[1],s_w_1);
AND_array_43 AND_array_43_c2({a_c[40:0],2'd0},p_prime[2],c_w_2);
AND_array_43 AND_array_43_s2({a_s[40:0],2'd0},p_prime[2],s_w_2);
AND_array_43 AND_array_43_c3({a_c[39:0],3'd0},p_prime[3],c_w_3);
AND_array_43 AND_array_43_s3({a_s[39:0],3'd0},p_prime[3],s_w_3);
AND_array_43 AND_array_43_c4({a_c[38:0],4'd0},p_prime[4],c_w_4);
AND_array_43 AND_array_43_s4({a_s[38:0],4'd0},p_prime[4],s_w_4);
AND_array_43 AND_array_43_c5({a_c[37:0],5'd0},p_prime[5],c_w_5);
AND_array_43 AND_array_43_s5({a_s[37:0],5'd0},p_prime[5],s_w_5);
AND_array_43 AND_array_43_c6({a_c[36:0],6'd0},p_prime[6],c_w_6);
AND_array_43 AND_array_43_s6({a_s[36:0],6'd0},p_prime[6],s_w_6);
AND_array_43 AND_array_43_c7({a_c[35:0],7'd0},p_prime[7],c_w_7);
AND_array_43 AND_array_43_s7({a_s[35:0],7'd0},p_prime[7],s_w_7);
AND_array_43 AND_array_43_c8({a_c[34:0],8'd0},p_prime[8],c_w_8);
AND_array_43 AND_array_43_s8({a_s[34:0],8'd0},p_prime[8],s_w_8);
AND_array_43 AND_array_43_c9({a_c[33:0],9'd0},p_prime[9],c_w_9);
AND_array_43 AND_array_43_s9({a_s[33:0],9'd0},p_prime[9],s_w_9);
AND_array_43 AND_array_43_c10({a_c[32:0],10'd0},p_prime[10],c_w_10);
AND_array_43 AND_array_43_s10({a_s[32:0],10'd0},p_prime[10],s_w_10);
AND_array_43 AND_array_43_c11({a_c[31:0],11'd0},p_prime[11],c_w_11);
AND_array_43 AND_array_43_s11({a_s[31:0],11'd0},p_prime[11],s_w_11);
AND_array_43 AND_array_43_c12({a_c[30:0],12'd0},p_prime[12],c_w_12);
AND_array_43 AND_array_43_s12({a_s[30:0],12'd0},p_prime[12],s_w_12);
AND_array_43 AND_array_43_c13({a_c[29:0],13'd0},p_prime[13],c_w_13);
AND_array_43 AND_array_43_s13({a_s[29:0],13'd0},p_prime[13],s_w_13);
AND_array_43 AND_array_43_c14({a_c[28:0],14'd0},p_prime[14],c_w_14);
AND_array_43 AND_array_43_s14({a_s[28:0],14'd0},p_prime[14],s_w_14);
AND_array_43 AND_array_43_c15({a_c[27:0],15'd0},p_prime[15],c_w_15);
AND_array_43 AND_array_43_s15({a_s[27:0],15'd0},p_prime[15],s_w_15);
AND_array_43 AND_array_43_c16({a_c[26:0],16'd0},p_prime[16],c_w_16);
AND_array_43 AND_array_43_s16({a_s[26:0],16'd0},p_prime[16],s_w_16);
AND_array_43 AND_array_43_c17({a_c[25:0],17'd0},p_prime[17],c_w_17);
AND_array_43 AND_array_43_s17({a_s[25:0],17'd0},p_prime[17],s_w_17);
AND_array_43 AND_array_43_c18({a_c[24:0],18'd0},p_prime[18],c_w_18);
AND_array_43 AND_array_43_s18({a_s[24:0],18'd0},p_prime[18],s_w_18);
AND_array_43 AND_array_43_c19({a_c[23:0],19'd0},p_prime[19],c_w_19);
AND_array_43 AND_array_43_s19({a_s[23:0],19'd0},p_prime[19],s_w_19);
AND_array_43 AND_array_43_c20({a_c[22:0],20'd0},p_prime[20],c_w_20);
AND_array_43 AND_array_43_s20({a_s[22:0],20'd0},p_prime[20],s_w_20);
AND_array_43 AND_array_43_c21({a_c[21:0],21'd0},p_prime[21],c_w_21);
AND_array_43 AND_array_43_s21({a_s[21:0],21'd0},p_prime[21],s_w_21);
AND_array_43 AND_array_43_c22({a_c[20:0],22'd0},p_prime[22],c_w_22);
AND_array_43 AND_array_43_s22({a_s[20:0],22'd0},p_prime[22],s_w_22);
AND_array_43 AND_array_43_c23({a_c[19:0],23'd0},p_prime[23],c_w_23);
AND_array_43 AND_array_43_s23({a_s[19:0],23'd0},p_prime[23],s_w_23);
AND_array_43 AND_array_43_c24({a_c[18:0],24'd0},p_prime[24],c_w_24);
AND_array_43 AND_array_43_s24({a_s[18:0],24'd0},p_prime[24],s_w_24);
AND_array_43 AND_array_43_c25({a_c[17:0],25'd0},p_prime[25],c_w_25);
AND_array_43 AND_array_43_s25({a_s[17:0],25'd0},p_prime[25],s_w_25);
AND_array_43 AND_array_43_c26({a_c[16:0],26'd0},p_prime[26],c_w_26);
AND_array_43 AND_array_43_s26({a_s[16:0],26'd0},p_prime[26],s_w_26);
AND_array_43 AND_array_43_c27({a_c[15:0],27'd0},p_prime[27],c_w_27);
AND_array_43 AND_array_43_s27({a_s[15:0],27'd0},p_prime[27],s_w_27);
AND_array_43 AND_array_43_c28({a_c[14:0],28'd0},p_prime[28],c_w_28);
AND_array_43 AND_array_43_s28({a_s[14:0],28'd0},p_prime[28],s_w_28);
AND_array_43 AND_array_43_c29({a_c[13:0],29'd0},p_prime[29],c_w_29);
AND_array_43 AND_array_43_s29({a_s[13:0],29'd0},p_prime[29],s_w_29);
AND_array_43 AND_array_43_c30({a_c[12:0],30'd0},p_prime[30],c_w_30);
AND_array_43 AND_array_43_s30({a_s[12:0],30'd0},p_prime[30],s_w_30);
AND_array_43 AND_array_43_c31({a_c[11:0],31'd0},p_prime[31],c_w_31);
AND_array_43 AND_array_43_s31({a_s[11:0],31'd0},p_prime[31],s_w_31);
AND_array_43 AND_array_43_c32({a_c[10:0],32'd0},p_prime[32],c_w_32);
AND_array_43 AND_array_43_s32({a_s[10:0],32'd0},p_prime[32],s_w_32);
AND_array_43 AND_array_43_c33({a_c[9:0],33'd0},p_prime[33],c_w_33);
AND_array_43 AND_array_43_s33({a_s[9:0],33'd0},p_prime[33],s_w_33);
AND_array_43 AND_array_43_c34({a_c[8:0],34'd0},p_prime[34],c_w_34);
AND_array_43 AND_array_43_s34({a_s[8:0],34'd0},p_prime[34],s_w_34);
AND_array_43 AND_array_43_c35({a_c[7:0],35'd0},p_prime[35],c_w_35);
AND_array_43 AND_array_43_s35({a_s[7:0],35'd0},p_prime[35],s_w_35);
AND_array_43 AND_array_43_c36({a_c[6:0],36'd0},p_prime[36],c_w_36);
AND_array_43 AND_array_43_s36({a_s[6:0],36'd0},p_prime[36],s_w_36);
AND_array_43 AND_array_43_c37({a_c[5:0],37'd0},p_prime[37],c_w_37);
AND_array_43 AND_array_43_s37({a_s[5:0],37'd0},p_prime[37],s_w_37);
AND_array_43 AND_array_43_c38({a_c[4:0],38'd0},p_prime[38],c_w_38);
AND_array_43 AND_array_43_s38({a_s[4:0],38'd0},p_prime[38],s_w_38);
AND_array_43 AND_array_43_c39({a_c[3:0],39'd0},p_prime[39],c_w_39);
AND_array_43 AND_array_43_s39({a_s[3:0],39'd0},p_prime[39],s_w_39);
AND_array_43 AND_array_43_c40({a_c[2:0],40'd0},p_prime[40],c_w_40);
AND_array_43 AND_array_43_s40({a_s[2:0],40'd0},p_prime[40],s_w_40);
AND_array_43 AND_array_43_c41({a_c[1:0],41'd0},p_prime[41],c_w_41);
AND_array_43 AND_array_43_s41({a_s[1:0],41'd0},p_prime[41],s_w_41);
AND_array_43 AND_array_43_c42({a_c[0:0],42'd0},p_prime[42],c_w_42);
AND_array_43 AND_array_43_s42({a_s[0:0],42'd0},p_prime[42],s_w_42);
    
assign b_c[42:0] = c_w_0;assign b_s[42:0] = s_w_0;
assign b_c[85:43] = c_w_1;assign b_s[85:43] = s_w_1;
assign b_c[128:86] = c_w_2;assign b_s[128:86] = s_w_2;
assign b_c[171:129] = c_w_3;assign b_s[171:129] = s_w_3;
assign b_c[214:172] = c_w_4;assign b_s[214:172] = s_w_4;
assign b_c[257:215] = c_w_5;assign b_s[257:215] = s_w_5;
assign b_c[300:258] = c_w_6;assign b_s[300:258] = s_w_6;
assign b_c[343:301] = c_w_7;assign b_s[343:301] = s_w_7;
assign b_c[386:344] = c_w_8;assign b_s[386:344] = s_w_8;
assign b_c[429:387] = c_w_9;assign b_s[429:387] = s_w_9;
assign b_c[472:430] = c_w_10;assign b_s[472:430] = s_w_10;
assign b_c[515:473] = c_w_11;assign b_s[515:473] = s_w_11;
assign b_c[558:516] = c_w_12;assign b_s[558:516] = s_w_12;
assign b_c[601:559] = c_w_13;assign b_s[601:559] = s_w_13;
assign b_c[644:602] = c_w_14;assign b_s[644:602] = s_w_14;
assign b_c[687:645] = c_w_15;assign b_s[687:645] = s_w_15;
assign b_c[730:688] = c_w_16;assign b_s[730:688] = s_w_16;
assign b_c[773:731] = c_w_17;assign b_s[773:731] = s_w_17;
assign b_c[816:774] = c_w_18;assign b_s[816:774] = s_w_18;
assign b_c[859:817] = c_w_19;assign b_s[859:817] = s_w_19;
assign b_c[902:860] = c_w_20;assign b_s[902:860] = s_w_20;
assign b_c[945:903] = c_w_21;assign b_s[945:903] = s_w_21;
assign b_c[988:946] = c_w_22;assign b_s[988:946] = s_w_22;
assign b_c[1031:989] = c_w_23;assign b_s[1031:989] = s_w_23;
assign b_c[1074:1032] = c_w_24;assign b_s[1074:1032] = s_w_24;
assign b_c[1117:1075] = c_w_25;assign b_s[1117:1075] = s_w_25;
assign b_c[1160:1118] = c_w_26;assign b_s[1160:1118] = s_w_26;
assign b_c[1203:1161] = c_w_27;assign b_s[1203:1161] = s_w_27;
assign b_c[1246:1204] = c_w_28;assign b_s[1246:1204] = s_w_28;
assign b_c[1289:1247] = c_w_29;assign b_s[1289:1247] = s_w_29;
assign b_c[1332:1290] = c_w_30;assign b_s[1332:1290] = s_w_30;
assign b_c[1375:1333] = c_w_31;assign b_s[1375:1333] = s_w_31;
assign b_c[1418:1376] = c_w_32;assign b_s[1418:1376] = s_w_32;
assign b_c[1461:1419] = c_w_33;assign b_s[1461:1419] = s_w_33;
assign b_c[1504:1462] = c_w_34;assign b_s[1504:1462] = s_w_34;
assign b_c[1547:1505] = c_w_35;assign b_s[1547:1505] = s_w_35;
assign b_c[1590:1548] = c_w_36;assign b_s[1590:1548] = s_w_36;
assign b_c[1633:1591] = c_w_37;assign b_s[1633:1591] = s_w_37;
assign b_c[1676:1634] = c_w_38;assign b_s[1676:1634] = s_w_38;
assign b_c[1719:1677] = c_w_39;assign b_s[1719:1677] = s_w_39;
assign b_c[1762:1720] = c_w_40;assign b_s[1762:1720] = s_w_40;
assign b_c[1805:1763] = c_w_41;assign b_s[1805:1763] = s_w_41;
assign b_c[1848:1806] = c_w_42;assign b_s[1848:1806] = s_w_42;
    
endmodule
    