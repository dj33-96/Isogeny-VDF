
module tb_4_iso_c_1506();

// Instruction list + effect:
/*
INS = 0 => Idle
INS = 1 => load input
INS = 2 => copy point rd to wr
INS = 3 => ADD
INS = 4 => SUB
INS = 5 => MUL
*/

reg clk,rst,get_output,data_en,ins_in;
wire [24-1:0] command_in;
reg [1506-1:0] din_1,din_2;
wire [1506-1:0] dout_1,dout_2;

reg [2:0] INS;
reg [7-1:0] rd_addr_1,rd_addr_2,wr_addr;

assign command_in = {INS,rd_addr_1,rd_addr_2,wr_addr};

wire [1506:0] p, calculated;
assign p = 1507'd1658539334852043956605014686969369842243820155059458240864380460354175875596746126442552006529285980003318752448184629099761975446397870870332614114924526019655624366944770281974501212314250998405682106067115619475132937730960746637418716661215852316737808364060021400361715167852784987427099666051667608448888314571788638487985846716927693574019769274326804364407638203115258648742883949562283207610572974523311143132532016594886767069744238342663307263;
assign calculated = (dout_1 + dout_2) % p;

wire [1506-1:0] x,z;//inputs
wire [1506-1:0] a,c,k1,k2,k3;//expected values

assign x = 1506'd940706300503281709855554913890461052139632021440893960843044572154501710007075923560090891594161561640555327597914143184810632733621040698095180777671697396567922467952258989868137440487306070421529612443442118761951018330734529996527053404562620107992031847886237842135094555234528562172726983127170853108419317392970192309174885112125304691730618936529983228422832446564425465780799213039184444161523251026993218759288219953527620155920296415270355175;
assign z = 1506'd612242396148598434486799786184741674417508768108009062352510425934148930985177095852531142164916640238348640109838023611753768331011788465977453770457014526026110708145667966514511288583025116710064481743298703213401248382965423952141059685844822097731389623578156025163412038802647435956351725731798369378465047961822199147767384444670405570437722454057189502255670765773895306607045324719378667166086720646121167292419043512143980672649925535370436085;
assign a = 1506'd275227671950079859646582086368814363894153200637395359178337690463517454154170491703638391639859105022146784401048868906882590799466275702897158648260500337624893146388018860817032217568179815107472377211721372227106398424004678509810376008809066660074049444921233924333020286897392224113591119903997603044461600883454108169916872860755148533792423093607506784011581252522605475499175549867217613527970361447226713514808045988613762585965912169044337802;
assign c = 1506'd1261155461947454011300267736388468063022232181216138077588521412715184536951805106536843170472130196359463195403130475485374879031935603902891601667347109508917363787258177358837516174013202347211420535856492649731758962343830506678908705358310742784431355184500023924326525384656812374992955605470832735987048072710865269506180123333216582025236092007643309044110410333836323585634131047886684981940518654511892544481420755136569030591286107531856218154;
assign k1 = 1506'd1539649505304839164296101196277002041699151911562988035801199524316123780866744278676539222231655627830222802795128678458793008834999421053669026250711916849992075241318187657985902706571535575136451745777611207308629368178148334155866127605317960711873959117122541996538228117534382623458733551909226852840214262687531686321964279983543850315950841196828377446508869192562614180394690347195967295170804495570907805531502384915181851645276638628530169421;
assign k2 = 1506'd328463904354683275368755127705719377722123253332884898490534146220352779021898827707559749429244921402206687488076119573056864402609252232117727007214682870541811759806591023353626151904280953711465130700143415548549769947769106044385993718717798010260642224308081816971682516431881126216375257395372483729954269431147993161407500667454899121292896482472793726167161680790530159173753888319805776995436530380872051466869176441383639483270370879899919090;
assign k3 = 1506'd1552948696651880144342354700075202726557140789548903023195554998088650640992253019412622033759078201878903967707752166796564401064632829164072634548128711922594033176097926956382648729070331187131594094186740821975352266713699953948668113090407442205723421471464393867298506594037175998129078708858969222486884365354792391456942269556795710262168341390587172730678503212338320772387844537758563111327609971673114386051707263465671600828570221950640791260;

cryptoprocessor_wrapper_1506 UUT(clk,rst,get_output,data_en,ins_in,command_in,din_1,din_2,dout_1,dout_2);

always #1 clk = ~clk;

initial begin
    clk = 0; rst = 0; data_en = 0; ins_in = 0; get_output = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd0,7'd0,7'd0,7'd0};
    @(posedge clk);
    rst = 1;get_output = 0;
    @(posedge clk);
    rst = 0;
    @(posedge clk);
    //Load x in addr 0
    data_en = 1; ins_in = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd1,7'd0,7'd0,7'd0};
    din_1 = x;
    din_2 = 0;
    @(posedge clk);
    //Load z in addr 1
    data_en = 1; ins_in = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd1,7'd0,7'd0,7'd1};
    din_1 = z;
    din_2 = 0;
    @(posedge clk);
    //Start the operations
    //addr5 = addr0 - addr1 | k2 = x - z
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd4,7'd0,7'd1,7'd5};
    @(posedge clk);
    //addr6 = addr0 + addr1 | k3 = x + z
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd3,7'd0,7'd1,7'd6};
    @(posedge clk);
    //addr4 = addr1 * addr1 | k1 = z ^ 2
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd1,7'd1,7'd4};
    @(posedge clk);
    //addr4 = addr4 + addr4 | k1 = k1 + k1
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd3,7'd4,7'd4,7'd4};
    @(posedge clk);
    //addr3 = addr4 * addr4 | c_iso = k1 ^ 2
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd4,7'd4,7'd3};
    @(posedge clk);
    //addr4 = addr4 + addr4 | k1 = k1 + k1
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd3,7'd4,7'd4,7'd4};
    @(posedge clk);
    //addr2 = addr0 * addr0 | a_iso = x ^ 2
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd0,7'd0,7'd2};
    @(posedge clk);
    //addr2 = addr2 + addr2 | a_iso = a_iso + a_iso
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd3,7'd2,7'd2,7'd2};
    @(posedge clk);
    //addr2 = addr2 * addr1 | a_iso = a_iso * a_iso
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd2,7'd2,7'd2};
    @(posedge clk);
    
    //Get output of addr = 2
    get_output = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd0,7'd2,7'd0,7'd0};
    @(posedge clk);
    if (a != calculated) begin
        $display("TEST for 4_iso_c: FAILED.");
        $display("Failed TEST: output = 0x%x,0x%x | a->4_iso_c = 0x%x, calculated = 0x%x",dout_1,dout_2,a,calculated);
        $display("Failed TEST: inputs: x,z = 0x%x,0x%x",x,z);
        $stop();
    end
    //Get output of addr = 3
    get_output = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd0,7'd3,7'd0,7'd0};
    @(posedge clk);
    if (c != calculated) begin
        $display("TEST for 4_iso_c: FAILED.");
        $display("Failed TEST: output = 0x%x,0x%x | c->4_iso_c = 0x%x, calculated = 0x%x",dout_1,dout_2,c,calculated);
        $display("Failed TEST: inputs: x,z = 0x%x,0x%x",x,z);
        $stop();
    end
    //Get output of addr = 4
    get_output = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd0,7'd4,7'd0,7'd0};
    @(posedge clk);
    if (k1%p != calculated%p) begin
        $display("TEST for 4_iso_c: FAILED.");
        $display("Failed TEST: output = 0x%x,0x%x | k1->4_iso_c = 0x%x, calculated = 0x%x",dout_1,dout_2,k1,calculated);
        $display("Failed TEST: inputs: x,z = 0x%x,0x%x",x,z);
        $stop();
    end
    //Get output of addr = 5
    get_output = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd0,7'd5,7'd0,7'd0};
    @(posedge clk);
    if (k2%p != calculated%p) begin
        $display("TEST for 4_iso_c: FAILED.");
        $display("Failed TEST: output = 0x%x,0x%x | k2->4_iso_c = 0x%x, calculated = 0x%x",dout_1,dout_2,k2,calculated);
        $display("Failed TEST: inputs: x,z = 0x%x,0x%x",x,z);
        $stop();
    end
    //Get output of addr = 6
    get_output = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd0,7'd6,7'd0,7'd0};
    @(posedge clk);
    if (k3%p != calculated%p) begin
        $display("TEST for 4_iso_c: FAILED.");
        $display("Failed TEST: output = 0x%x,0x%x | k3->4_iso_c = 0x%x, calculated = 0x%x",dout_1,dout_2,k3,calculated);
        $display("Failed TEST: inputs: x,z = 0x%x,0x%x",x,z);
        $stop();
    end
    @(posedge clk);
    
    $display("4-iso-c correct");
    $finish();
end

endmodule
    