

module csa_tree_40x80(
    input [3199:0] A, // lines are appended together
    output[79:0] B_0,
    output[79:0] B_1
);

wire [2159:0] tree_1;
wire [1439:0] tree_2;
wire [959:0] tree_3;
wire [639:0] tree_4;
wire [479:0] tree_5;
wire [319:0] tree_6;
wire [239:0] tree_7;
wire [159:0] tree_8;
// layer-1
csa_80 csau_80_i0(A[79:0],A[159:80],A[239:160],tree_1[79:0],tree_1[159:80]);
csa_80 csau_80_i1(A[319:240],A[399:320],A[479:400],tree_1[239:160],tree_1[319:240]);
csa_80 csau_80_i2(A[559:480],A[639:560],A[719:640],tree_1[399:320],tree_1[479:400]);
csa_80 csau_80_i3(A[799:720],A[879:800],A[959:880],tree_1[559:480],tree_1[639:560]);
csa_80 csau_80_i4(A[1039:960],A[1119:1040],A[1199:1120],tree_1[719:640],tree_1[799:720]);
csa_80 csau_80_i5(A[1279:1200],A[1359:1280],A[1439:1360],tree_1[879:800],tree_1[959:880]);
csa_80 csau_80_i6(A[1519:1440],A[1599:1520],A[1679:1600],tree_1[1039:960],tree_1[1119:1040]);
csa_80 csau_80_i7(A[1759:1680],A[1839:1760],A[1919:1840],tree_1[1199:1120],tree_1[1279:1200]);
csa_80 csau_80_i8(A[1999:1920],A[2079:2000],A[2159:2080],tree_1[1359:1280],tree_1[1439:1360]);
csa_80 csau_80_i9(A[2239:2160],A[2319:2240],A[2399:2320],tree_1[1519:1440],tree_1[1599:1520]);
csa_80 csau_80_i10(A[2479:2400],A[2559:2480],A[2639:2560],tree_1[1679:1600],tree_1[1759:1680]);
csa_80 csau_80_i11(A[2719:2640],A[2799:2720],A[2879:2800],tree_1[1839:1760],tree_1[1919:1840]);
csa_80 csau_80_i12(A[2959:2880],A[3039:2960],A[3119:3040],tree_1[1999:1920],tree_1[2079:2000]);
assign tree_1[2159:2080] = A[3199:3120];
// layer-2
csa_80 csau_80_i13(tree_1[79:0],tree_1[159:80],tree_1[239:160],tree_2[79:0],tree_2[159:80]);
csa_80 csau_80_i14(tree_1[319:240],tree_1[399:320],tree_1[479:400],tree_2[239:160],tree_2[319:240]);
csa_80 csau_80_i15(tree_1[559:480],tree_1[639:560],tree_1[719:640],tree_2[399:320],tree_2[479:400]);
csa_80 csau_80_i16(tree_1[799:720],tree_1[879:800],tree_1[959:880],tree_2[559:480],tree_2[639:560]);
csa_80 csau_80_i17(tree_1[1039:960],tree_1[1119:1040],tree_1[1199:1120],tree_2[719:640],tree_2[799:720]);
csa_80 csau_80_i18(tree_1[1279:1200],tree_1[1359:1280],tree_1[1439:1360],tree_2[879:800],tree_2[959:880]);
csa_80 csau_80_i19(tree_1[1519:1440],tree_1[1599:1520],tree_1[1679:1600],tree_2[1039:960],tree_2[1119:1040]);
csa_80 csau_80_i20(tree_1[1759:1680],tree_1[1839:1760],tree_1[1919:1840],tree_2[1199:1120],tree_2[1279:1200]);
csa_80 csau_80_i21(tree_1[1999:1920],tree_1[2079:2000],tree_1[2159:2080],tree_2[1359:1280],tree_2[1439:1360]);
// layer-3
csa_80 csau_80_i22(tree_2[79:0],tree_2[159:80],tree_2[239:160],tree_3[79:0],tree_3[159:80]);
csa_80 csau_80_i23(tree_2[319:240],tree_2[399:320],tree_2[479:400],tree_3[239:160],tree_3[319:240]);
csa_80 csau_80_i24(tree_2[559:480],tree_2[639:560],tree_2[719:640],tree_3[399:320],tree_3[479:400]);
csa_80 csau_80_i25(tree_2[799:720],tree_2[879:800],tree_2[959:880],tree_3[559:480],tree_3[639:560]);
csa_80 csau_80_i26(tree_2[1039:960],tree_2[1119:1040],tree_2[1199:1120],tree_3[719:640],tree_3[799:720]);
csa_80 csau_80_i27(tree_2[1279:1200],tree_2[1359:1280],tree_2[1439:1360],tree_3[879:800],tree_3[959:880]);
// layer-4
csa_80 csau_80_i28(tree_3[79:0],tree_3[159:80],tree_3[239:160],tree_4[79:0],tree_4[159:80]);
csa_80 csau_80_i29(tree_3[319:240],tree_3[399:320],tree_3[479:400],tree_4[239:160],tree_4[319:240]);
csa_80 csau_80_i30(tree_3[559:480],tree_3[639:560],tree_3[719:640],tree_4[399:320],tree_4[479:400]);
csa_80 csau_80_i31(tree_3[799:720],tree_3[879:800],tree_3[959:880],tree_4[559:480],tree_4[639:560]);
// layer-5
csa_80 csau_80_i32(tree_4[79:0],tree_4[159:80],tree_4[239:160],tree_5[79:0],tree_5[159:80]);
csa_80 csau_80_i33(tree_4[319:240],tree_4[399:320],tree_4[479:400],tree_5[239:160],tree_5[319:240]);
assign tree_5[399:320] = tree_4[559:480];
assign tree_5[479:400] = tree_4[639:560];
// layer-6
csa_80 csau_80_i34(tree_5[79:0],tree_5[159:80],tree_5[239:160],tree_6[79:0],tree_6[159:80]);
csa_80 csau_80_i35(tree_5[319:240],tree_5[399:320],tree_5[479:400],tree_6[239:160],tree_6[319:240]);
// layer-7
csa_80 csau_80_i36(tree_6[79:0],tree_6[159:80],tree_6[239:160],tree_7[79:0],tree_7[159:80]);
assign tree_7[239:160] = tree_6[319:240];
// layer-8
csa_80 csau_80_i37(tree_7[79:0],tree_7[159:80],tree_7[239:160],tree_8[79:0],tree_8[159:80]);

// final assignment
assign B_0 = tree_8[79:0];
assign B_1 = tree_8[159:80];

endmodule
