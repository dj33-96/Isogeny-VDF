
module AND_matrix_89x89(
    input [88:0] a,
    input [88:0] b,
    output [15841:0] c // lines are appended together
);
    
wire [88:0] c_w_0;
wire [88:0] c_w_1;
wire [88:0] c_w_2;
wire [88:0] c_w_3;
wire [88:0] c_w_4;
wire [88:0] c_w_5;
wire [88:0] c_w_6;
wire [88:0] c_w_7;
wire [88:0] c_w_8;
wire [88:0] c_w_9;
wire [88:0] c_w_10;
wire [88:0] c_w_11;
wire [88:0] c_w_12;
wire [88:0] c_w_13;
wire [88:0] c_w_14;
wire [88:0] c_w_15;
wire [88:0] c_w_16;
wire [88:0] c_w_17;
wire [88:0] c_w_18;
wire [88:0] c_w_19;
wire [88:0] c_w_20;
wire [88:0] c_w_21;
wire [88:0] c_w_22;
wire [88:0] c_w_23;
wire [88:0] c_w_24;
wire [88:0] c_w_25;
wire [88:0] c_w_26;
wire [88:0] c_w_27;
wire [88:0] c_w_28;
wire [88:0] c_w_29;
wire [88:0] c_w_30;
wire [88:0] c_w_31;
wire [88:0] c_w_32;
wire [88:0] c_w_33;
wire [88:0] c_w_34;
wire [88:0] c_w_35;
wire [88:0] c_w_36;
wire [88:0] c_w_37;
wire [88:0] c_w_38;
wire [88:0] c_w_39;
wire [88:0] c_w_40;
wire [88:0] c_w_41;
wire [88:0] c_w_42;
wire [88:0] c_w_43;
wire [88:0] c_w_44;
wire [88:0] c_w_45;
wire [88:0] c_w_46;
wire [88:0] c_w_47;
wire [88:0] c_w_48;
wire [88:0] c_w_49;
wire [88:0] c_w_50;
wire [88:0] c_w_51;
wire [88:0] c_w_52;
wire [88:0] c_w_53;
wire [88:0] c_w_54;
wire [88:0] c_w_55;
wire [88:0] c_w_56;
wire [88:0] c_w_57;
wire [88:0] c_w_58;
wire [88:0] c_w_59;
wire [88:0] c_w_60;
wire [88:0] c_w_61;
wire [88:0] c_w_62;
wire [88:0] c_w_63;
wire [88:0] c_w_64;
wire [88:0] c_w_65;
wire [88:0] c_w_66;
wire [88:0] c_w_67;
wire [88:0] c_w_68;
wire [88:0] c_w_69;
wire [88:0] c_w_70;
wire [88:0] c_w_71;
wire [88:0] c_w_72;
wire [88:0] c_w_73;
wire [88:0] c_w_74;
wire [88:0] c_w_75;
wire [88:0] c_w_76;
wire [88:0] c_w_77;
wire [88:0] c_w_78;
wire [88:0] c_w_79;
wire [88:0] c_w_80;
wire [88:0] c_w_81;
wire [88:0] c_w_82;
wire [88:0] c_w_83;
wire [88:0] c_w_84;
wire [88:0] c_w_85;
wire [88:0] c_w_86;
wire [88:0] c_w_87;
wire [88:0] c_w_88;
    
AND_array_89 AND_array_89_i0(a,b[0],c_w_0);
AND_array_89 AND_array_89_i1(a,b[1],c_w_1);
AND_array_89 AND_array_89_i2(a,b[2],c_w_2);
AND_array_89 AND_array_89_i3(a,b[3],c_w_3);
AND_array_89 AND_array_89_i4(a,b[4],c_w_4);
AND_array_89 AND_array_89_i5(a,b[5],c_w_5);
AND_array_89 AND_array_89_i6(a,b[6],c_w_6);
AND_array_89 AND_array_89_i7(a,b[7],c_w_7);
AND_array_89 AND_array_89_i8(a,b[8],c_w_8);
AND_array_89 AND_array_89_i9(a,b[9],c_w_9);
AND_array_89 AND_array_89_i10(a,b[10],c_w_10);
AND_array_89 AND_array_89_i11(a,b[11],c_w_11);
AND_array_89 AND_array_89_i12(a,b[12],c_w_12);
AND_array_89 AND_array_89_i13(a,b[13],c_w_13);
AND_array_89 AND_array_89_i14(a,b[14],c_w_14);
AND_array_89 AND_array_89_i15(a,b[15],c_w_15);
AND_array_89 AND_array_89_i16(a,b[16],c_w_16);
AND_array_89 AND_array_89_i17(a,b[17],c_w_17);
AND_array_89 AND_array_89_i18(a,b[18],c_w_18);
AND_array_89 AND_array_89_i19(a,b[19],c_w_19);
AND_array_89 AND_array_89_i20(a,b[20],c_w_20);
AND_array_89 AND_array_89_i21(a,b[21],c_w_21);
AND_array_89 AND_array_89_i22(a,b[22],c_w_22);
AND_array_89 AND_array_89_i23(a,b[23],c_w_23);
AND_array_89 AND_array_89_i24(a,b[24],c_w_24);
AND_array_89 AND_array_89_i25(a,b[25],c_w_25);
AND_array_89 AND_array_89_i26(a,b[26],c_w_26);
AND_array_89 AND_array_89_i27(a,b[27],c_w_27);
AND_array_89 AND_array_89_i28(a,b[28],c_w_28);
AND_array_89 AND_array_89_i29(a,b[29],c_w_29);
AND_array_89 AND_array_89_i30(a,b[30],c_w_30);
AND_array_89 AND_array_89_i31(a,b[31],c_w_31);
AND_array_89 AND_array_89_i32(a,b[32],c_w_32);
AND_array_89 AND_array_89_i33(a,b[33],c_w_33);
AND_array_89 AND_array_89_i34(a,b[34],c_w_34);
AND_array_89 AND_array_89_i35(a,b[35],c_w_35);
AND_array_89 AND_array_89_i36(a,b[36],c_w_36);
AND_array_89 AND_array_89_i37(a,b[37],c_w_37);
AND_array_89 AND_array_89_i38(a,b[38],c_w_38);
AND_array_89 AND_array_89_i39(a,b[39],c_w_39);
AND_array_89 AND_array_89_i40(a,b[40],c_w_40);
AND_array_89 AND_array_89_i41(a,b[41],c_w_41);
AND_array_89 AND_array_89_i42(a,b[42],c_w_42);
AND_array_89 AND_array_89_i43(a,b[43],c_w_43);
AND_array_89 AND_array_89_i44(a,b[44],c_w_44);
AND_array_89 AND_array_89_i45(a,b[45],c_w_45);
AND_array_89 AND_array_89_i46(a,b[46],c_w_46);
AND_array_89 AND_array_89_i47(a,b[47],c_w_47);
AND_array_89 AND_array_89_i48(a,b[48],c_w_48);
AND_array_89 AND_array_89_i49(a,b[49],c_w_49);
AND_array_89 AND_array_89_i50(a,b[50],c_w_50);
AND_array_89 AND_array_89_i51(a,b[51],c_w_51);
AND_array_89 AND_array_89_i52(a,b[52],c_w_52);
AND_array_89 AND_array_89_i53(a,b[53],c_w_53);
AND_array_89 AND_array_89_i54(a,b[54],c_w_54);
AND_array_89 AND_array_89_i55(a,b[55],c_w_55);
AND_array_89 AND_array_89_i56(a,b[56],c_w_56);
AND_array_89 AND_array_89_i57(a,b[57],c_w_57);
AND_array_89 AND_array_89_i58(a,b[58],c_w_58);
AND_array_89 AND_array_89_i59(a,b[59],c_w_59);
AND_array_89 AND_array_89_i60(a,b[60],c_w_60);
AND_array_89 AND_array_89_i61(a,b[61],c_w_61);
AND_array_89 AND_array_89_i62(a,b[62],c_w_62);
AND_array_89 AND_array_89_i63(a,b[63],c_w_63);
AND_array_89 AND_array_89_i64(a,b[64],c_w_64);
AND_array_89 AND_array_89_i65(a,b[65],c_w_65);
AND_array_89 AND_array_89_i66(a,b[66],c_w_66);
AND_array_89 AND_array_89_i67(a,b[67],c_w_67);
AND_array_89 AND_array_89_i68(a,b[68],c_w_68);
AND_array_89 AND_array_89_i69(a,b[69],c_w_69);
AND_array_89 AND_array_89_i70(a,b[70],c_w_70);
AND_array_89 AND_array_89_i71(a,b[71],c_w_71);
AND_array_89 AND_array_89_i72(a,b[72],c_w_72);
AND_array_89 AND_array_89_i73(a,b[73],c_w_73);
AND_array_89 AND_array_89_i74(a,b[74],c_w_74);
AND_array_89 AND_array_89_i75(a,b[75],c_w_75);
AND_array_89 AND_array_89_i76(a,b[76],c_w_76);
AND_array_89 AND_array_89_i77(a,b[77],c_w_77);
AND_array_89 AND_array_89_i78(a,b[78],c_w_78);
AND_array_89 AND_array_89_i79(a,b[79],c_w_79);
AND_array_89 AND_array_89_i80(a,b[80],c_w_80);
AND_array_89 AND_array_89_i81(a,b[81],c_w_81);
AND_array_89 AND_array_89_i82(a,b[82],c_w_82);
AND_array_89 AND_array_89_i83(a,b[83],c_w_83);
AND_array_89 AND_array_89_i84(a,b[84],c_w_84);
AND_array_89 AND_array_89_i85(a,b[85],c_w_85);
AND_array_89 AND_array_89_i86(a,b[86],c_w_86);
AND_array_89 AND_array_89_i87(a,b[87],c_w_87);
AND_array_89 AND_array_89_i88(a,b[88],c_w_88);
    
assign c[177:0] = {89'b0,c_w_0};
assign c[355:178] = {88'b0,c_w_1,1'b0};
assign c[533:356] = {87'b0,c_w_2,2'b0};
assign c[711:534] = {86'b0,c_w_3,3'b0};
assign c[889:712] = {85'b0,c_w_4,4'b0};
assign c[1067:890] = {84'b0,c_w_5,5'b0};
assign c[1245:1068] = {83'b0,c_w_6,6'b0};
assign c[1423:1246] = {82'b0,c_w_7,7'b0};
assign c[1601:1424] = {81'b0,c_w_8,8'b0};
assign c[1779:1602] = {80'b0,c_w_9,9'b0};
assign c[1957:1780] = {79'b0,c_w_10,10'b0};
assign c[2135:1958] = {78'b0,c_w_11,11'b0};
assign c[2313:2136] = {77'b0,c_w_12,12'b0};
assign c[2491:2314] = {76'b0,c_w_13,13'b0};
assign c[2669:2492] = {75'b0,c_w_14,14'b0};
assign c[2847:2670] = {74'b0,c_w_15,15'b0};
assign c[3025:2848] = {73'b0,c_w_16,16'b0};
assign c[3203:3026] = {72'b0,c_w_17,17'b0};
assign c[3381:3204] = {71'b0,c_w_18,18'b0};
assign c[3559:3382] = {70'b0,c_w_19,19'b0};
assign c[3737:3560] = {69'b0,c_w_20,20'b0};
assign c[3915:3738] = {68'b0,c_w_21,21'b0};
assign c[4093:3916] = {67'b0,c_w_22,22'b0};
assign c[4271:4094] = {66'b0,c_w_23,23'b0};
assign c[4449:4272] = {65'b0,c_w_24,24'b0};
assign c[4627:4450] = {64'b0,c_w_25,25'b0};
assign c[4805:4628] = {63'b0,c_w_26,26'b0};
assign c[4983:4806] = {62'b0,c_w_27,27'b0};
assign c[5161:4984] = {61'b0,c_w_28,28'b0};
assign c[5339:5162] = {60'b0,c_w_29,29'b0};
assign c[5517:5340] = {59'b0,c_w_30,30'b0};
assign c[5695:5518] = {58'b0,c_w_31,31'b0};
assign c[5873:5696] = {57'b0,c_w_32,32'b0};
assign c[6051:5874] = {56'b0,c_w_33,33'b0};
assign c[6229:6052] = {55'b0,c_w_34,34'b0};
assign c[6407:6230] = {54'b0,c_w_35,35'b0};
assign c[6585:6408] = {53'b0,c_w_36,36'b0};
assign c[6763:6586] = {52'b0,c_w_37,37'b0};
assign c[6941:6764] = {51'b0,c_w_38,38'b0};
assign c[7119:6942] = {50'b0,c_w_39,39'b0};
assign c[7297:7120] = {49'b0,c_w_40,40'b0};
assign c[7475:7298] = {48'b0,c_w_41,41'b0};
assign c[7653:7476] = {47'b0,c_w_42,42'b0};
assign c[7831:7654] = {46'b0,c_w_43,43'b0};
assign c[8009:7832] = {45'b0,c_w_44,44'b0};
assign c[8187:8010] = {44'b0,c_w_45,45'b0};
assign c[8365:8188] = {43'b0,c_w_46,46'b0};
assign c[8543:8366] = {42'b0,c_w_47,47'b0};
assign c[8721:8544] = {41'b0,c_w_48,48'b0};
assign c[8899:8722] = {40'b0,c_w_49,49'b0};
assign c[9077:8900] = {39'b0,c_w_50,50'b0};
assign c[9255:9078] = {38'b0,c_w_51,51'b0};
assign c[9433:9256] = {37'b0,c_w_52,52'b0};
assign c[9611:9434] = {36'b0,c_w_53,53'b0};
assign c[9789:9612] = {35'b0,c_w_54,54'b0};
assign c[9967:9790] = {34'b0,c_w_55,55'b0};
assign c[10145:9968] = {33'b0,c_w_56,56'b0};
assign c[10323:10146] = {32'b0,c_w_57,57'b0};
assign c[10501:10324] = {31'b0,c_w_58,58'b0};
assign c[10679:10502] = {30'b0,c_w_59,59'b0};
assign c[10857:10680] = {29'b0,c_w_60,60'b0};
assign c[11035:10858] = {28'b0,c_w_61,61'b0};
assign c[11213:11036] = {27'b0,c_w_62,62'b0};
assign c[11391:11214] = {26'b0,c_w_63,63'b0};
assign c[11569:11392] = {25'b0,c_w_64,64'b0};
assign c[11747:11570] = {24'b0,c_w_65,65'b0};
assign c[11925:11748] = {23'b0,c_w_66,66'b0};
assign c[12103:11926] = {22'b0,c_w_67,67'b0};
assign c[12281:12104] = {21'b0,c_w_68,68'b0};
assign c[12459:12282] = {20'b0,c_w_69,69'b0};
assign c[12637:12460] = {19'b0,c_w_70,70'b0};
assign c[12815:12638] = {18'b0,c_w_71,71'b0};
assign c[12993:12816] = {17'b0,c_w_72,72'b0};
assign c[13171:12994] = {16'b0,c_w_73,73'b0};
assign c[13349:13172] = {15'b0,c_w_74,74'b0};
assign c[13527:13350] = {14'b0,c_w_75,75'b0};
assign c[13705:13528] = {13'b0,c_w_76,76'b0};
assign c[13883:13706] = {12'b0,c_w_77,77'b0};
assign c[14061:13884] = {11'b0,c_w_78,78'b0};
assign c[14239:14062] = {10'b0,c_w_79,79'b0};
assign c[14417:14240] = {9'b0,c_w_80,80'b0};
assign c[14595:14418] = {8'b0,c_w_81,81'b0};
assign c[14773:14596] = {7'b0,c_w_82,82'b0};
assign c[14951:14774] = {6'b0,c_w_83,83'b0};
assign c[15129:14952] = {5'b0,c_w_84,84'b0};
assign c[15307:15130] = {4'b0,c_w_85,85'b0};
assign c[15485:15308] = {3'b0,c_w_86,86'b0};
assign c[15663:15486] = {2'b0,c_w_87,87'b0};
assign c[15841:15664] = {1'b0,c_w_88,88'b0};
    
endmodule
    