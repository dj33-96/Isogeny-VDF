
module xor_1506_array(
    input [1505:0] in0,in1,
    output [1505:0] out0
);

assign out0 = in0 ^ in1;

endmodule
    