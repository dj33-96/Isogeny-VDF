
module add_1506_lut(
    input [2:0] M,
    output reg [1505:0] corr_add
);

always @(*) begin
    case(M)
    3'd0: corr_add = 1506'h0;
    3'd1: corr_add = 1506'h20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    3'd2: corr_add = 1506'h10b6cad46b6070b7ed381d9cea88c74ea092c836403f32b6eb2ac931cabd9bd2a300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
    3'd3: corr_add = 1506'h16d95a8d6c0e16fda703b39d5118e9d4125906c807e656dd6559263957b37a54600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002;
    3'd4: corr_add = 1506'h216d95a8d6c0e16fda703b39d5118e9d4125906c807e656dd6559263957b37a54600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002;
    3'd5: corr_add = 1506'h1224607d42215227c7a858d6bf9a55ebe1b858a2c0bd9824c1805b956038d377e900000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003;
    3'd6: corr_add = 1506'h2db2b51ad81c2dfb4e07673aa231d3a824b20d900fccadbacab24c72af66f4a8c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004;
    3'd7: corr_add = 1506'h22db2b51ad81c2dfb4e07673aa231d3a824b20d900fccadbacab24c72af66f4a8c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004;
    default: corr_add = 0;
    endcase
end

endmodule
    