
module csa_3018 (
    input [3017:0] x,y,z,
    output[3017:0] c,s 
);

wire dummy;

assign c[0] = 1'b0;
    
assign {c[1],s[0]} = (x[0]+y[0]+z[0]);
assign {c[2],s[1]} = (x[1]+y[1]+z[1]);
assign {c[3],s[2]} = (x[2]+y[2]+z[2]);
assign {c[4],s[3]} = (x[3]+y[3]+z[3]);
assign {c[5],s[4]} = (x[4]+y[4]+z[4]);
assign {c[6],s[5]} = (x[5]+y[5]+z[5]);
assign {c[7],s[6]} = (x[6]+y[6]+z[6]);
assign {c[8],s[7]} = (x[7]+y[7]+z[7]);
assign {c[9],s[8]} = (x[8]+y[8]+z[8]);
assign {c[10],s[9]} = (x[9]+y[9]+z[9]);
assign {c[11],s[10]} = (x[10]+y[10]+z[10]);
assign {c[12],s[11]} = (x[11]+y[11]+z[11]);
assign {c[13],s[12]} = (x[12]+y[12]+z[12]);
assign {c[14],s[13]} = (x[13]+y[13]+z[13]);
assign {c[15],s[14]} = (x[14]+y[14]+z[14]);
assign {c[16],s[15]} = (x[15]+y[15]+z[15]);
assign {c[17],s[16]} = (x[16]+y[16]+z[16]);
assign {c[18],s[17]} = (x[17]+y[17]+z[17]);
assign {c[19],s[18]} = (x[18]+y[18]+z[18]);
assign {c[20],s[19]} = (x[19]+y[19]+z[19]);
assign {c[21],s[20]} = (x[20]+y[20]+z[20]);
assign {c[22],s[21]} = (x[21]+y[21]+z[21]);
assign {c[23],s[22]} = (x[22]+y[22]+z[22]);
assign {c[24],s[23]} = (x[23]+y[23]+z[23]);
assign {c[25],s[24]} = (x[24]+y[24]+z[24]);
assign {c[26],s[25]} = (x[25]+y[25]+z[25]);
assign {c[27],s[26]} = (x[26]+y[26]+z[26]);
assign {c[28],s[27]} = (x[27]+y[27]+z[27]);
assign {c[29],s[28]} = (x[28]+y[28]+z[28]);
assign {c[30],s[29]} = (x[29]+y[29]+z[29]);
assign {c[31],s[30]} = (x[30]+y[30]+z[30]);
assign {c[32],s[31]} = (x[31]+y[31]+z[31]);
assign {c[33],s[32]} = (x[32]+y[32]+z[32]);
assign {c[34],s[33]} = (x[33]+y[33]+z[33]);
assign {c[35],s[34]} = (x[34]+y[34]+z[34]);
assign {c[36],s[35]} = (x[35]+y[35]+z[35]);
assign {c[37],s[36]} = (x[36]+y[36]+z[36]);
assign {c[38],s[37]} = (x[37]+y[37]+z[37]);
assign {c[39],s[38]} = (x[38]+y[38]+z[38]);
assign {c[40],s[39]} = (x[39]+y[39]+z[39]);
assign {c[41],s[40]} = (x[40]+y[40]+z[40]);
assign {c[42],s[41]} = (x[41]+y[41]+z[41]);
assign {c[43],s[42]} = (x[42]+y[42]+z[42]);
assign {c[44],s[43]} = (x[43]+y[43]+z[43]);
assign {c[45],s[44]} = (x[44]+y[44]+z[44]);
assign {c[46],s[45]} = (x[45]+y[45]+z[45]);
assign {c[47],s[46]} = (x[46]+y[46]+z[46]);
assign {c[48],s[47]} = (x[47]+y[47]+z[47]);
assign {c[49],s[48]} = (x[48]+y[48]+z[48]);
assign {c[50],s[49]} = (x[49]+y[49]+z[49]);
assign {c[51],s[50]} = (x[50]+y[50]+z[50]);
assign {c[52],s[51]} = (x[51]+y[51]+z[51]);
assign {c[53],s[52]} = (x[52]+y[52]+z[52]);
assign {c[54],s[53]} = (x[53]+y[53]+z[53]);
assign {c[55],s[54]} = (x[54]+y[54]+z[54]);
assign {c[56],s[55]} = (x[55]+y[55]+z[55]);
assign {c[57],s[56]} = (x[56]+y[56]+z[56]);
assign {c[58],s[57]} = (x[57]+y[57]+z[57]);
assign {c[59],s[58]} = (x[58]+y[58]+z[58]);
assign {c[60],s[59]} = (x[59]+y[59]+z[59]);
assign {c[61],s[60]} = (x[60]+y[60]+z[60]);
assign {c[62],s[61]} = (x[61]+y[61]+z[61]);
assign {c[63],s[62]} = (x[62]+y[62]+z[62]);
assign {c[64],s[63]} = (x[63]+y[63]+z[63]);
assign {c[65],s[64]} = (x[64]+y[64]+z[64]);
assign {c[66],s[65]} = (x[65]+y[65]+z[65]);
assign {c[67],s[66]} = (x[66]+y[66]+z[66]);
assign {c[68],s[67]} = (x[67]+y[67]+z[67]);
assign {c[69],s[68]} = (x[68]+y[68]+z[68]);
assign {c[70],s[69]} = (x[69]+y[69]+z[69]);
assign {c[71],s[70]} = (x[70]+y[70]+z[70]);
assign {c[72],s[71]} = (x[71]+y[71]+z[71]);
assign {c[73],s[72]} = (x[72]+y[72]+z[72]);
assign {c[74],s[73]} = (x[73]+y[73]+z[73]);
assign {c[75],s[74]} = (x[74]+y[74]+z[74]);
assign {c[76],s[75]} = (x[75]+y[75]+z[75]);
assign {c[77],s[76]} = (x[76]+y[76]+z[76]);
assign {c[78],s[77]} = (x[77]+y[77]+z[77]);
assign {c[79],s[78]} = (x[78]+y[78]+z[78]);
assign {c[80],s[79]} = (x[79]+y[79]+z[79]);
assign {c[81],s[80]} = (x[80]+y[80]+z[80]);
assign {c[82],s[81]} = (x[81]+y[81]+z[81]);
assign {c[83],s[82]} = (x[82]+y[82]+z[82]);
assign {c[84],s[83]} = (x[83]+y[83]+z[83]);
assign {c[85],s[84]} = (x[84]+y[84]+z[84]);
assign {c[86],s[85]} = (x[85]+y[85]+z[85]);
assign {c[87],s[86]} = (x[86]+y[86]+z[86]);
assign {c[88],s[87]} = (x[87]+y[87]+z[87]);
assign {c[89],s[88]} = (x[88]+y[88]+z[88]);
assign {c[90],s[89]} = (x[89]+y[89]+z[89]);
assign {c[91],s[90]} = (x[90]+y[90]+z[90]);
assign {c[92],s[91]} = (x[91]+y[91]+z[91]);
assign {c[93],s[92]} = (x[92]+y[92]+z[92]);
assign {c[94],s[93]} = (x[93]+y[93]+z[93]);
assign {c[95],s[94]} = (x[94]+y[94]+z[94]);
assign {c[96],s[95]} = (x[95]+y[95]+z[95]);
assign {c[97],s[96]} = (x[96]+y[96]+z[96]);
assign {c[98],s[97]} = (x[97]+y[97]+z[97]);
assign {c[99],s[98]} = (x[98]+y[98]+z[98]);
assign {c[100],s[99]} = (x[99]+y[99]+z[99]);
assign {c[101],s[100]} = (x[100]+y[100]+z[100]);
assign {c[102],s[101]} = (x[101]+y[101]+z[101]);
assign {c[103],s[102]} = (x[102]+y[102]+z[102]);
assign {c[104],s[103]} = (x[103]+y[103]+z[103]);
assign {c[105],s[104]} = (x[104]+y[104]+z[104]);
assign {c[106],s[105]} = (x[105]+y[105]+z[105]);
assign {c[107],s[106]} = (x[106]+y[106]+z[106]);
assign {c[108],s[107]} = (x[107]+y[107]+z[107]);
assign {c[109],s[108]} = (x[108]+y[108]+z[108]);
assign {c[110],s[109]} = (x[109]+y[109]+z[109]);
assign {c[111],s[110]} = (x[110]+y[110]+z[110]);
assign {c[112],s[111]} = (x[111]+y[111]+z[111]);
assign {c[113],s[112]} = (x[112]+y[112]+z[112]);
assign {c[114],s[113]} = (x[113]+y[113]+z[113]);
assign {c[115],s[114]} = (x[114]+y[114]+z[114]);
assign {c[116],s[115]} = (x[115]+y[115]+z[115]);
assign {c[117],s[116]} = (x[116]+y[116]+z[116]);
assign {c[118],s[117]} = (x[117]+y[117]+z[117]);
assign {c[119],s[118]} = (x[118]+y[118]+z[118]);
assign {c[120],s[119]} = (x[119]+y[119]+z[119]);
assign {c[121],s[120]} = (x[120]+y[120]+z[120]);
assign {c[122],s[121]} = (x[121]+y[121]+z[121]);
assign {c[123],s[122]} = (x[122]+y[122]+z[122]);
assign {c[124],s[123]} = (x[123]+y[123]+z[123]);
assign {c[125],s[124]} = (x[124]+y[124]+z[124]);
assign {c[126],s[125]} = (x[125]+y[125]+z[125]);
assign {c[127],s[126]} = (x[126]+y[126]+z[126]);
assign {c[128],s[127]} = (x[127]+y[127]+z[127]);
assign {c[129],s[128]} = (x[128]+y[128]+z[128]);
assign {c[130],s[129]} = (x[129]+y[129]+z[129]);
assign {c[131],s[130]} = (x[130]+y[130]+z[130]);
assign {c[132],s[131]} = (x[131]+y[131]+z[131]);
assign {c[133],s[132]} = (x[132]+y[132]+z[132]);
assign {c[134],s[133]} = (x[133]+y[133]+z[133]);
assign {c[135],s[134]} = (x[134]+y[134]+z[134]);
assign {c[136],s[135]} = (x[135]+y[135]+z[135]);
assign {c[137],s[136]} = (x[136]+y[136]+z[136]);
assign {c[138],s[137]} = (x[137]+y[137]+z[137]);
assign {c[139],s[138]} = (x[138]+y[138]+z[138]);
assign {c[140],s[139]} = (x[139]+y[139]+z[139]);
assign {c[141],s[140]} = (x[140]+y[140]+z[140]);
assign {c[142],s[141]} = (x[141]+y[141]+z[141]);
assign {c[143],s[142]} = (x[142]+y[142]+z[142]);
assign {c[144],s[143]} = (x[143]+y[143]+z[143]);
assign {c[145],s[144]} = (x[144]+y[144]+z[144]);
assign {c[146],s[145]} = (x[145]+y[145]+z[145]);
assign {c[147],s[146]} = (x[146]+y[146]+z[146]);
assign {c[148],s[147]} = (x[147]+y[147]+z[147]);
assign {c[149],s[148]} = (x[148]+y[148]+z[148]);
assign {c[150],s[149]} = (x[149]+y[149]+z[149]);
assign {c[151],s[150]} = (x[150]+y[150]+z[150]);
assign {c[152],s[151]} = (x[151]+y[151]+z[151]);
assign {c[153],s[152]} = (x[152]+y[152]+z[152]);
assign {c[154],s[153]} = (x[153]+y[153]+z[153]);
assign {c[155],s[154]} = (x[154]+y[154]+z[154]);
assign {c[156],s[155]} = (x[155]+y[155]+z[155]);
assign {c[157],s[156]} = (x[156]+y[156]+z[156]);
assign {c[158],s[157]} = (x[157]+y[157]+z[157]);
assign {c[159],s[158]} = (x[158]+y[158]+z[158]);
assign {c[160],s[159]} = (x[159]+y[159]+z[159]);
assign {c[161],s[160]} = (x[160]+y[160]+z[160]);
assign {c[162],s[161]} = (x[161]+y[161]+z[161]);
assign {c[163],s[162]} = (x[162]+y[162]+z[162]);
assign {c[164],s[163]} = (x[163]+y[163]+z[163]);
assign {c[165],s[164]} = (x[164]+y[164]+z[164]);
assign {c[166],s[165]} = (x[165]+y[165]+z[165]);
assign {c[167],s[166]} = (x[166]+y[166]+z[166]);
assign {c[168],s[167]} = (x[167]+y[167]+z[167]);
assign {c[169],s[168]} = (x[168]+y[168]+z[168]);
assign {c[170],s[169]} = (x[169]+y[169]+z[169]);
assign {c[171],s[170]} = (x[170]+y[170]+z[170]);
assign {c[172],s[171]} = (x[171]+y[171]+z[171]);
assign {c[173],s[172]} = (x[172]+y[172]+z[172]);
assign {c[174],s[173]} = (x[173]+y[173]+z[173]);
assign {c[175],s[174]} = (x[174]+y[174]+z[174]);
assign {c[176],s[175]} = (x[175]+y[175]+z[175]);
assign {c[177],s[176]} = (x[176]+y[176]+z[176]);
assign {c[178],s[177]} = (x[177]+y[177]+z[177]);
assign {c[179],s[178]} = (x[178]+y[178]+z[178]);
assign {c[180],s[179]} = (x[179]+y[179]+z[179]);
assign {c[181],s[180]} = (x[180]+y[180]+z[180]);
assign {c[182],s[181]} = (x[181]+y[181]+z[181]);
assign {c[183],s[182]} = (x[182]+y[182]+z[182]);
assign {c[184],s[183]} = (x[183]+y[183]+z[183]);
assign {c[185],s[184]} = (x[184]+y[184]+z[184]);
assign {c[186],s[185]} = (x[185]+y[185]+z[185]);
assign {c[187],s[186]} = (x[186]+y[186]+z[186]);
assign {c[188],s[187]} = (x[187]+y[187]+z[187]);
assign {c[189],s[188]} = (x[188]+y[188]+z[188]);
assign {c[190],s[189]} = (x[189]+y[189]+z[189]);
assign {c[191],s[190]} = (x[190]+y[190]+z[190]);
assign {c[192],s[191]} = (x[191]+y[191]+z[191]);
assign {c[193],s[192]} = (x[192]+y[192]+z[192]);
assign {c[194],s[193]} = (x[193]+y[193]+z[193]);
assign {c[195],s[194]} = (x[194]+y[194]+z[194]);
assign {c[196],s[195]} = (x[195]+y[195]+z[195]);
assign {c[197],s[196]} = (x[196]+y[196]+z[196]);
assign {c[198],s[197]} = (x[197]+y[197]+z[197]);
assign {c[199],s[198]} = (x[198]+y[198]+z[198]);
assign {c[200],s[199]} = (x[199]+y[199]+z[199]);
assign {c[201],s[200]} = (x[200]+y[200]+z[200]);
assign {c[202],s[201]} = (x[201]+y[201]+z[201]);
assign {c[203],s[202]} = (x[202]+y[202]+z[202]);
assign {c[204],s[203]} = (x[203]+y[203]+z[203]);
assign {c[205],s[204]} = (x[204]+y[204]+z[204]);
assign {c[206],s[205]} = (x[205]+y[205]+z[205]);
assign {c[207],s[206]} = (x[206]+y[206]+z[206]);
assign {c[208],s[207]} = (x[207]+y[207]+z[207]);
assign {c[209],s[208]} = (x[208]+y[208]+z[208]);
assign {c[210],s[209]} = (x[209]+y[209]+z[209]);
assign {c[211],s[210]} = (x[210]+y[210]+z[210]);
assign {c[212],s[211]} = (x[211]+y[211]+z[211]);
assign {c[213],s[212]} = (x[212]+y[212]+z[212]);
assign {c[214],s[213]} = (x[213]+y[213]+z[213]);
assign {c[215],s[214]} = (x[214]+y[214]+z[214]);
assign {c[216],s[215]} = (x[215]+y[215]+z[215]);
assign {c[217],s[216]} = (x[216]+y[216]+z[216]);
assign {c[218],s[217]} = (x[217]+y[217]+z[217]);
assign {c[219],s[218]} = (x[218]+y[218]+z[218]);
assign {c[220],s[219]} = (x[219]+y[219]+z[219]);
assign {c[221],s[220]} = (x[220]+y[220]+z[220]);
assign {c[222],s[221]} = (x[221]+y[221]+z[221]);
assign {c[223],s[222]} = (x[222]+y[222]+z[222]);
assign {c[224],s[223]} = (x[223]+y[223]+z[223]);
assign {c[225],s[224]} = (x[224]+y[224]+z[224]);
assign {c[226],s[225]} = (x[225]+y[225]+z[225]);
assign {c[227],s[226]} = (x[226]+y[226]+z[226]);
assign {c[228],s[227]} = (x[227]+y[227]+z[227]);
assign {c[229],s[228]} = (x[228]+y[228]+z[228]);
assign {c[230],s[229]} = (x[229]+y[229]+z[229]);
assign {c[231],s[230]} = (x[230]+y[230]+z[230]);
assign {c[232],s[231]} = (x[231]+y[231]+z[231]);
assign {c[233],s[232]} = (x[232]+y[232]+z[232]);
assign {c[234],s[233]} = (x[233]+y[233]+z[233]);
assign {c[235],s[234]} = (x[234]+y[234]+z[234]);
assign {c[236],s[235]} = (x[235]+y[235]+z[235]);
assign {c[237],s[236]} = (x[236]+y[236]+z[236]);
assign {c[238],s[237]} = (x[237]+y[237]+z[237]);
assign {c[239],s[238]} = (x[238]+y[238]+z[238]);
assign {c[240],s[239]} = (x[239]+y[239]+z[239]);
assign {c[241],s[240]} = (x[240]+y[240]+z[240]);
assign {c[242],s[241]} = (x[241]+y[241]+z[241]);
assign {c[243],s[242]} = (x[242]+y[242]+z[242]);
assign {c[244],s[243]} = (x[243]+y[243]+z[243]);
assign {c[245],s[244]} = (x[244]+y[244]+z[244]);
assign {c[246],s[245]} = (x[245]+y[245]+z[245]);
assign {c[247],s[246]} = (x[246]+y[246]+z[246]);
assign {c[248],s[247]} = (x[247]+y[247]+z[247]);
assign {c[249],s[248]} = (x[248]+y[248]+z[248]);
assign {c[250],s[249]} = (x[249]+y[249]+z[249]);
assign {c[251],s[250]} = (x[250]+y[250]+z[250]);
assign {c[252],s[251]} = (x[251]+y[251]+z[251]);
assign {c[253],s[252]} = (x[252]+y[252]+z[252]);
assign {c[254],s[253]} = (x[253]+y[253]+z[253]);
assign {c[255],s[254]} = (x[254]+y[254]+z[254]);
assign {c[256],s[255]} = (x[255]+y[255]+z[255]);
assign {c[257],s[256]} = (x[256]+y[256]+z[256]);
assign {c[258],s[257]} = (x[257]+y[257]+z[257]);
assign {c[259],s[258]} = (x[258]+y[258]+z[258]);
assign {c[260],s[259]} = (x[259]+y[259]+z[259]);
assign {c[261],s[260]} = (x[260]+y[260]+z[260]);
assign {c[262],s[261]} = (x[261]+y[261]+z[261]);
assign {c[263],s[262]} = (x[262]+y[262]+z[262]);
assign {c[264],s[263]} = (x[263]+y[263]+z[263]);
assign {c[265],s[264]} = (x[264]+y[264]+z[264]);
assign {c[266],s[265]} = (x[265]+y[265]+z[265]);
assign {c[267],s[266]} = (x[266]+y[266]+z[266]);
assign {c[268],s[267]} = (x[267]+y[267]+z[267]);
assign {c[269],s[268]} = (x[268]+y[268]+z[268]);
assign {c[270],s[269]} = (x[269]+y[269]+z[269]);
assign {c[271],s[270]} = (x[270]+y[270]+z[270]);
assign {c[272],s[271]} = (x[271]+y[271]+z[271]);
assign {c[273],s[272]} = (x[272]+y[272]+z[272]);
assign {c[274],s[273]} = (x[273]+y[273]+z[273]);
assign {c[275],s[274]} = (x[274]+y[274]+z[274]);
assign {c[276],s[275]} = (x[275]+y[275]+z[275]);
assign {c[277],s[276]} = (x[276]+y[276]+z[276]);
assign {c[278],s[277]} = (x[277]+y[277]+z[277]);
assign {c[279],s[278]} = (x[278]+y[278]+z[278]);
assign {c[280],s[279]} = (x[279]+y[279]+z[279]);
assign {c[281],s[280]} = (x[280]+y[280]+z[280]);
assign {c[282],s[281]} = (x[281]+y[281]+z[281]);
assign {c[283],s[282]} = (x[282]+y[282]+z[282]);
assign {c[284],s[283]} = (x[283]+y[283]+z[283]);
assign {c[285],s[284]} = (x[284]+y[284]+z[284]);
assign {c[286],s[285]} = (x[285]+y[285]+z[285]);
assign {c[287],s[286]} = (x[286]+y[286]+z[286]);
assign {c[288],s[287]} = (x[287]+y[287]+z[287]);
assign {c[289],s[288]} = (x[288]+y[288]+z[288]);
assign {c[290],s[289]} = (x[289]+y[289]+z[289]);
assign {c[291],s[290]} = (x[290]+y[290]+z[290]);
assign {c[292],s[291]} = (x[291]+y[291]+z[291]);
assign {c[293],s[292]} = (x[292]+y[292]+z[292]);
assign {c[294],s[293]} = (x[293]+y[293]+z[293]);
assign {c[295],s[294]} = (x[294]+y[294]+z[294]);
assign {c[296],s[295]} = (x[295]+y[295]+z[295]);
assign {c[297],s[296]} = (x[296]+y[296]+z[296]);
assign {c[298],s[297]} = (x[297]+y[297]+z[297]);
assign {c[299],s[298]} = (x[298]+y[298]+z[298]);
assign {c[300],s[299]} = (x[299]+y[299]+z[299]);
assign {c[301],s[300]} = (x[300]+y[300]+z[300]);
assign {c[302],s[301]} = (x[301]+y[301]+z[301]);
assign {c[303],s[302]} = (x[302]+y[302]+z[302]);
assign {c[304],s[303]} = (x[303]+y[303]+z[303]);
assign {c[305],s[304]} = (x[304]+y[304]+z[304]);
assign {c[306],s[305]} = (x[305]+y[305]+z[305]);
assign {c[307],s[306]} = (x[306]+y[306]+z[306]);
assign {c[308],s[307]} = (x[307]+y[307]+z[307]);
assign {c[309],s[308]} = (x[308]+y[308]+z[308]);
assign {c[310],s[309]} = (x[309]+y[309]+z[309]);
assign {c[311],s[310]} = (x[310]+y[310]+z[310]);
assign {c[312],s[311]} = (x[311]+y[311]+z[311]);
assign {c[313],s[312]} = (x[312]+y[312]+z[312]);
assign {c[314],s[313]} = (x[313]+y[313]+z[313]);
assign {c[315],s[314]} = (x[314]+y[314]+z[314]);
assign {c[316],s[315]} = (x[315]+y[315]+z[315]);
assign {c[317],s[316]} = (x[316]+y[316]+z[316]);
assign {c[318],s[317]} = (x[317]+y[317]+z[317]);
assign {c[319],s[318]} = (x[318]+y[318]+z[318]);
assign {c[320],s[319]} = (x[319]+y[319]+z[319]);
assign {c[321],s[320]} = (x[320]+y[320]+z[320]);
assign {c[322],s[321]} = (x[321]+y[321]+z[321]);
assign {c[323],s[322]} = (x[322]+y[322]+z[322]);
assign {c[324],s[323]} = (x[323]+y[323]+z[323]);
assign {c[325],s[324]} = (x[324]+y[324]+z[324]);
assign {c[326],s[325]} = (x[325]+y[325]+z[325]);
assign {c[327],s[326]} = (x[326]+y[326]+z[326]);
assign {c[328],s[327]} = (x[327]+y[327]+z[327]);
assign {c[329],s[328]} = (x[328]+y[328]+z[328]);
assign {c[330],s[329]} = (x[329]+y[329]+z[329]);
assign {c[331],s[330]} = (x[330]+y[330]+z[330]);
assign {c[332],s[331]} = (x[331]+y[331]+z[331]);
assign {c[333],s[332]} = (x[332]+y[332]+z[332]);
assign {c[334],s[333]} = (x[333]+y[333]+z[333]);
assign {c[335],s[334]} = (x[334]+y[334]+z[334]);
assign {c[336],s[335]} = (x[335]+y[335]+z[335]);
assign {c[337],s[336]} = (x[336]+y[336]+z[336]);
assign {c[338],s[337]} = (x[337]+y[337]+z[337]);
assign {c[339],s[338]} = (x[338]+y[338]+z[338]);
assign {c[340],s[339]} = (x[339]+y[339]+z[339]);
assign {c[341],s[340]} = (x[340]+y[340]+z[340]);
assign {c[342],s[341]} = (x[341]+y[341]+z[341]);
assign {c[343],s[342]} = (x[342]+y[342]+z[342]);
assign {c[344],s[343]} = (x[343]+y[343]+z[343]);
assign {c[345],s[344]} = (x[344]+y[344]+z[344]);
assign {c[346],s[345]} = (x[345]+y[345]+z[345]);
assign {c[347],s[346]} = (x[346]+y[346]+z[346]);
assign {c[348],s[347]} = (x[347]+y[347]+z[347]);
assign {c[349],s[348]} = (x[348]+y[348]+z[348]);
assign {c[350],s[349]} = (x[349]+y[349]+z[349]);
assign {c[351],s[350]} = (x[350]+y[350]+z[350]);
assign {c[352],s[351]} = (x[351]+y[351]+z[351]);
assign {c[353],s[352]} = (x[352]+y[352]+z[352]);
assign {c[354],s[353]} = (x[353]+y[353]+z[353]);
assign {c[355],s[354]} = (x[354]+y[354]+z[354]);
assign {c[356],s[355]} = (x[355]+y[355]+z[355]);
assign {c[357],s[356]} = (x[356]+y[356]+z[356]);
assign {c[358],s[357]} = (x[357]+y[357]+z[357]);
assign {c[359],s[358]} = (x[358]+y[358]+z[358]);
assign {c[360],s[359]} = (x[359]+y[359]+z[359]);
assign {c[361],s[360]} = (x[360]+y[360]+z[360]);
assign {c[362],s[361]} = (x[361]+y[361]+z[361]);
assign {c[363],s[362]} = (x[362]+y[362]+z[362]);
assign {c[364],s[363]} = (x[363]+y[363]+z[363]);
assign {c[365],s[364]} = (x[364]+y[364]+z[364]);
assign {c[366],s[365]} = (x[365]+y[365]+z[365]);
assign {c[367],s[366]} = (x[366]+y[366]+z[366]);
assign {c[368],s[367]} = (x[367]+y[367]+z[367]);
assign {c[369],s[368]} = (x[368]+y[368]+z[368]);
assign {c[370],s[369]} = (x[369]+y[369]+z[369]);
assign {c[371],s[370]} = (x[370]+y[370]+z[370]);
assign {c[372],s[371]} = (x[371]+y[371]+z[371]);
assign {c[373],s[372]} = (x[372]+y[372]+z[372]);
assign {c[374],s[373]} = (x[373]+y[373]+z[373]);
assign {c[375],s[374]} = (x[374]+y[374]+z[374]);
assign {c[376],s[375]} = (x[375]+y[375]+z[375]);
assign {c[377],s[376]} = (x[376]+y[376]+z[376]);
assign {c[378],s[377]} = (x[377]+y[377]+z[377]);
assign {c[379],s[378]} = (x[378]+y[378]+z[378]);
assign {c[380],s[379]} = (x[379]+y[379]+z[379]);
assign {c[381],s[380]} = (x[380]+y[380]+z[380]);
assign {c[382],s[381]} = (x[381]+y[381]+z[381]);
assign {c[383],s[382]} = (x[382]+y[382]+z[382]);
assign {c[384],s[383]} = (x[383]+y[383]+z[383]);
assign {c[385],s[384]} = (x[384]+y[384]+z[384]);
assign {c[386],s[385]} = (x[385]+y[385]+z[385]);
assign {c[387],s[386]} = (x[386]+y[386]+z[386]);
assign {c[388],s[387]} = (x[387]+y[387]+z[387]);
assign {c[389],s[388]} = (x[388]+y[388]+z[388]);
assign {c[390],s[389]} = (x[389]+y[389]+z[389]);
assign {c[391],s[390]} = (x[390]+y[390]+z[390]);
assign {c[392],s[391]} = (x[391]+y[391]+z[391]);
assign {c[393],s[392]} = (x[392]+y[392]+z[392]);
assign {c[394],s[393]} = (x[393]+y[393]+z[393]);
assign {c[395],s[394]} = (x[394]+y[394]+z[394]);
assign {c[396],s[395]} = (x[395]+y[395]+z[395]);
assign {c[397],s[396]} = (x[396]+y[396]+z[396]);
assign {c[398],s[397]} = (x[397]+y[397]+z[397]);
assign {c[399],s[398]} = (x[398]+y[398]+z[398]);
assign {c[400],s[399]} = (x[399]+y[399]+z[399]);
assign {c[401],s[400]} = (x[400]+y[400]+z[400]);
assign {c[402],s[401]} = (x[401]+y[401]+z[401]);
assign {c[403],s[402]} = (x[402]+y[402]+z[402]);
assign {c[404],s[403]} = (x[403]+y[403]+z[403]);
assign {c[405],s[404]} = (x[404]+y[404]+z[404]);
assign {c[406],s[405]} = (x[405]+y[405]+z[405]);
assign {c[407],s[406]} = (x[406]+y[406]+z[406]);
assign {c[408],s[407]} = (x[407]+y[407]+z[407]);
assign {c[409],s[408]} = (x[408]+y[408]+z[408]);
assign {c[410],s[409]} = (x[409]+y[409]+z[409]);
assign {c[411],s[410]} = (x[410]+y[410]+z[410]);
assign {c[412],s[411]} = (x[411]+y[411]+z[411]);
assign {c[413],s[412]} = (x[412]+y[412]+z[412]);
assign {c[414],s[413]} = (x[413]+y[413]+z[413]);
assign {c[415],s[414]} = (x[414]+y[414]+z[414]);
assign {c[416],s[415]} = (x[415]+y[415]+z[415]);
assign {c[417],s[416]} = (x[416]+y[416]+z[416]);
assign {c[418],s[417]} = (x[417]+y[417]+z[417]);
assign {c[419],s[418]} = (x[418]+y[418]+z[418]);
assign {c[420],s[419]} = (x[419]+y[419]+z[419]);
assign {c[421],s[420]} = (x[420]+y[420]+z[420]);
assign {c[422],s[421]} = (x[421]+y[421]+z[421]);
assign {c[423],s[422]} = (x[422]+y[422]+z[422]);
assign {c[424],s[423]} = (x[423]+y[423]+z[423]);
assign {c[425],s[424]} = (x[424]+y[424]+z[424]);
assign {c[426],s[425]} = (x[425]+y[425]+z[425]);
assign {c[427],s[426]} = (x[426]+y[426]+z[426]);
assign {c[428],s[427]} = (x[427]+y[427]+z[427]);
assign {c[429],s[428]} = (x[428]+y[428]+z[428]);
assign {c[430],s[429]} = (x[429]+y[429]+z[429]);
assign {c[431],s[430]} = (x[430]+y[430]+z[430]);
assign {c[432],s[431]} = (x[431]+y[431]+z[431]);
assign {c[433],s[432]} = (x[432]+y[432]+z[432]);
assign {c[434],s[433]} = (x[433]+y[433]+z[433]);
assign {c[435],s[434]} = (x[434]+y[434]+z[434]);
assign {c[436],s[435]} = (x[435]+y[435]+z[435]);
assign {c[437],s[436]} = (x[436]+y[436]+z[436]);
assign {c[438],s[437]} = (x[437]+y[437]+z[437]);
assign {c[439],s[438]} = (x[438]+y[438]+z[438]);
assign {c[440],s[439]} = (x[439]+y[439]+z[439]);
assign {c[441],s[440]} = (x[440]+y[440]+z[440]);
assign {c[442],s[441]} = (x[441]+y[441]+z[441]);
assign {c[443],s[442]} = (x[442]+y[442]+z[442]);
assign {c[444],s[443]} = (x[443]+y[443]+z[443]);
assign {c[445],s[444]} = (x[444]+y[444]+z[444]);
assign {c[446],s[445]} = (x[445]+y[445]+z[445]);
assign {c[447],s[446]} = (x[446]+y[446]+z[446]);
assign {c[448],s[447]} = (x[447]+y[447]+z[447]);
assign {c[449],s[448]} = (x[448]+y[448]+z[448]);
assign {c[450],s[449]} = (x[449]+y[449]+z[449]);
assign {c[451],s[450]} = (x[450]+y[450]+z[450]);
assign {c[452],s[451]} = (x[451]+y[451]+z[451]);
assign {c[453],s[452]} = (x[452]+y[452]+z[452]);
assign {c[454],s[453]} = (x[453]+y[453]+z[453]);
assign {c[455],s[454]} = (x[454]+y[454]+z[454]);
assign {c[456],s[455]} = (x[455]+y[455]+z[455]);
assign {c[457],s[456]} = (x[456]+y[456]+z[456]);
assign {c[458],s[457]} = (x[457]+y[457]+z[457]);
assign {c[459],s[458]} = (x[458]+y[458]+z[458]);
assign {c[460],s[459]} = (x[459]+y[459]+z[459]);
assign {c[461],s[460]} = (x[460]+y[460]+z[460]);
assign {c[462],s[461]} = (x[461]+y[461]+z[461]);
assign {c[463],s[462]} = (x[462]+y[462]+z[462]);
assign {c[464],s[463]} = (x[463]+y[463]+z[463]);
assign {c[465],s[464]} = (x[464]+y[464]+z[464]);
assign {c[466],s[465]} = (x[465]+y[465]+z[465]);
assign {c[467],s[466]} = (x[466]+y[466]+z[466]);
assign {c[468],s[467]} = (x[467]+y[467]+z[467]);
assign {c[469],s[468]} = (x[468]+y[468]+z[468]);
assign {c[470],s[469]} = (x[469]+y[469]+z[469]);
assign {c[471],s[470]} = (x[470]+y[470]+z[470]);
assign {c[472],s[471]} = (x[471]+y[471]+z[471]);
assign {c[473],s[472]} = (x[472]+y[472]+z[472]);
assign {c[474],s[473]} = (x[473]+y[473]+z[473]);
assign {c[475],s[474]} = (x[474]+y[474]+z[474]);
assign {c[476],s[475]} = (x[475]+y[475]+z[475]);
assign {c[477],s[476]} = (x[476]+y[476]+z[476]);
assign {c[478],s[477]} = (x[477]+y[477]+z[477]);
assign {c[479],s[478]} = (x[478]+y[478]+z[478]);
assign {c[480],s[479]} = (x[479]+y[479]+z[479]);
assign {c[481],s[480]} = (x[480]+y[480]+z[480]);
assign {c[482],s[481]} = (x[481]+y[481]+z[481]);
assign {c[483],s[482]} = (x[482]+y[482]+z[482]);
assign {c[484],s[483]} = (x[483]+y[483]+z[483]);
assign {c[485],s[484]} = (x[484]+y[484]+z[484]);
assign {c[486],s[485]} = (x[485]+y[485]+z[485]);
assign {c[487],s[486]} = (x[486]+y[486]+z[486]);
assign {c[488],s[487]} = (x[487]+y[487]+z[487]);
assign {c[489],s[488]} = (x[488]+y[488]+z[488]);
assign {c[490],s[489]} = (x[489]+y[489]+z[489]);
assign {c[491],s[490]} = (x[490]+y[490]+z[490]);
assign {c[492],s[491]} = (x[491]+y[491]+z[491]);
assign {c[493],s[492]} = (x[492]+y[492]+z[492]);
assign {c[494],s[493]} = (x[493]+y[493]+z[493]);
assign {c[495],s[494]} = (x[494]+y[494]+z[494]);
assign {c[496],s[495]} = (x[495]+y[495]+z[495]);
assign {c[497],s[496]} = (x[496]+y[496]+z[496]);
assign {c[498],s[497]} = (x[497]+y[497]+z[497]);
assign {c[499],s[498]} = (x[498]+y[498]+z[498]);
assign {c[500],s[499]} = (x[499]+y[499]+z[499]);
assign {c[501],s[500]} = (x[500]+y[500]+z[500]);
assign {c[502],s[501]} = (x[501]+y[501]+z[501]);
assign {c[503],s[502]} = (x[502]+y[502]+z[502]);
assign {c[504],s[503]} = (x[503]+y[503]+z[503]);
assign {c[505],s[504]} = (x[504]+y[504]+z[504]);
assign {c[506],s[505]} = (x[505]+y[505]+z[505]);
assign {c[507],s[506]} = (x[506]+y[506]+z[506]);
assign {c[508],s[507]} = (x[507]+y[507]+z[507]);
assign {c[509],s[508]} = (x[508]+y[508]+z[508]);
assign {c[510],s[509]} = (x[509]+y[509]+z[509]);
assign {c[511],s[510]} = (x[510]+y[510]+z[510]);
assign {c[512],s[511]} = (x[511]+y[511]+z[511]);
assign {c[513],s[512]} = (x[512]+y[512]+z[512]);
assign {c[514],s[513]} = (x[513]+y[513]+z[513]);
assign {c[515],s[514]} = (x[514]+y[514]+z[514]);
assign {c[516],s[515]} = (x[515]+y[515]+z[515]);
assign {c[517],s[516]} = (x[516]+y[516]+z[516]);
assign {c[518],s[517]} = (x[517]+y[517]+z[517]);
assign {c[519],s[518]} = (x[518]+y[518]+z[518]);
assign {c[520],s[519]} = (x[519]+y[519]+z[519]);
assign {c[521],s[520]} = (x[520]+y[520]+z[520]);
assign {c[522],s[521]} = (x[521]+y[521]+z[521]);
assign {c[523],s[522]} = (x[522]+y[522]+z[522]);
assign {c[524],s[523]} = (x[523]+y[523]+z[523]);
assign {c[525],s[524]} = (x[524]+y[524]+z[524]);
assign {c[526],s[525]} = (x[525]+y[525]+z[525]);
assign {c[527],s[526]} = (x[526]+y[526]+z[526]);
assign {c[528],s[527]} = (x[527]+y[527]+z[527]);
assign {c[529],s[528]} = (x[528]+y[528]+z[528]);
assign {c[530],s[529]} = (x[529]+y[529]+z[529]);
assign {c[531],s[530]} = (x[530]+y[530]+z[530]);
assign {c[532],s[531]} = (x[531]+y[531]+z[531]);
assign {c[533],s[532]} = (x[532]+y[532]+z[532]);
assign {c[534],s[533]} = (x[533]+y[533]+z[533]);
assign {c[535],s[534]} = (x[534]+y[534]+z[534]);
assign {c[536],s[535]} = (x[535]+y[535]+z[535]);
assign {c[537],s[536]} = (x[536]+y[536]+z[536]);
assign {c[538],s[537]} = (x[537]+y[537]+z[537]);
assign {c[539],s[538]} = (x[538]+y[538]+z[538]);
assign {c[540],s[539]} = (x[539]+y[539]+z[539]);
assign {c[541],s[540]} = (x[540]+y[540]+z[540]);
assign {c[542],s[541]} = (x[541]+y[541]+z[541]);
assign {c[543],s[542]} = (x[542]+y[542]+z[542]);
assign {c[544],s[543]} = (x[543]+y[543]+z[543]);
assign {c[545],s[544]} = (x[544]+y[544]+z[544]);
assign {c[546],s[545]} = (x[545]+y[545]+z[545]);
assign {c[547],s[546]} = (x[546]+y[546]+z[546]);
assign {c[548],s[547]} = (x[547]+y[547]+z[547]);
assign {c[549],s[548]} = (x[548]+y[548]+z[548]);
assign {c[550],s[549]} = (x[549]+y[549]+z[549]);
assign {c[551],s[550]} = (x[550]+y[550]+z[550]);
assign {c[552],s[551]} = (x[551]+y[551]+z[551]);
assign {c[553],s[552]} = (x[552]+y[552]+z[552]);
assign {c[554],s[553]} = (x[553]+y[553]+z[553]);
assign {c[555],s[554]} = (x[554]+y[554]+z[554]);
assign {c[556],s[555]} = (x[555]+y[555]+z[555]);
assign {c[557],s[556]} = (x[556]+y[556]+z[556]);
assign {c[558],s[557]} = (x[557]+y[557]+z[557]);
assign {c[559],s[558]} = (x[558]+y[558]+z[558]);
assign {c[560],s[559]} = (x[559]+y[559]+z[559]);
assign {c[561],s[560]} = (x[560]+y[560]+z[560]);
assign {c[562],s[561]} = (x[561]+y[561]+z[561]);
assign {c[563],s[562]} = (x[562]+y[562]+z[562]);
assign {c[564],s[563]} = (x[563]+y[563]+z[563]);
assign {c[565],s[564]} = (x[564]+y[564]+z[564]);
assign {c[566],s[565]} = (x[565]+y[565]+z[565]);
assign {c[567],s[566]} = (x[566]+y[566]+z[566]);
assign {c[568],s[567]} = (x[567]+y[567]+z[567]);
assign {c[569],s[568]} = (x[568]+y[568]+z[568]);
assign {c[570],s[569]} = (x[569]+y[569]+z[569]);
assign {c[571],s[570]} = (x[570]+y[570]+z[570]);
assign {c[572],s[571]} = (x[571]+y[571]+z[571]);
assign {c[573],s[572]} = (x[572]+y[572]+z[572]);
assign {c[574],s[573]} = (x[573]+y[573]+z[573]);
assign {c[575],s[574]} = (x[574]+y[574]+z[574]);
assign {c[576],s[575]} = (x[575]+y[575]+z[575]);
assign {c[577],s[576]} = (x[576]+y[576]+z[576]);
assign {c[578],s[577]} = (x[577]+y[577]+z[577]);
assign {c[579],s[578]} = (x[578]+y[578]+z[578]);
assign {c[580],s[579]} = (x[579]+y[579]+z[579]);
assign {c[581],s[580]} = (x[580]+y[580]+z[580]);
assign {c[582],s[581]} = (x[581]+y[581]+z[581]);
assign {c[583],s[582]} = (x[582]+y[582]+z[582]);
assign {c[584],s[583]} = (x[583]+y[583]+z[583]);
assign {c[585],s[584]} = (x[584]+y[584]+z[584]);
assign {c[586],s[585]} = (x[585]+y[585]+z[585]);
assign {c[587],s[586]} = (x[586]+y[586]+z[586]);
assign {c[588],s[587]} = (x[587]+y[587]+z[587]);
assign {c[589],s[588]} = (x[588]+y[588]+z[588]);
assign {c[590],s[589]} = (x[589]+y[589]+z[589]);
assign {c[591],s[590]} = (x[590]+y[590]+z[590]);
assign {c[592],s[591]} = (x[591]+y[591]+z[591]);
assign {c[593],s[592]} = (x[592]+y[592]+z[592]);
assign {c[594],s[593]} = (x[593]+y[593]+z[593]);
assign {c[595],s[594]} = (x[594]+y[594]+z[594]);
assign {c[596],s[595]} = (x[595]+y[595]+z[595]);
assign {c[597],s[596]} = (x[596]+y[596]+z[596]);
assign {c[598],s[597]} = (x[597]+y[597]+z[597]);
assign {c[599],s[598]} = (x[598]+y[598]+z[598]);
assign {c[600],s[599]} = (x[599]+y[599]+z[599]);
assign {c[601],s[600]} = (x[600]+y[600]+z[600]);
assign {c[602],s[601]} = (x[601]+y[601]+z[601]);
assign {c[603],s[602]} = (x[602]+y[602]+z[602]);
assign {c[604],s[603]} = (x[603]+y[603]+z[603]);
assign {c[605],s[604]} = (x[604]+y[604]+z[604]);
assign {c[606],s[605]} = (x[605]+y[605]+z[605]);
assign {c[607],s[606]} = (x[606]+y[606]+z[606]);
assign {c[608],s[607]} = (x[607]+y[607]+z[607]);
assign {c[609],s[608]} = (x[608]+y[608]+z[608]);
assign {c[610],s[609]} = (x[609]+y[609]+z[609]);
assign {c[611],s[610]} = (x[610]+y[610]+z[610]);
assign {c[612],s[611]} = (x[611]+y[611]+z[611]);
assign {c[613],s[612]} = (x[612]+y[612]+z[612]);
assign {c[614],s[613]} = (x[613]+y[613]+z[613]);
assign {c[615],s[614]} = (x[614]+y[614]+z[614]);
assign {c[616],s[615]} = (x[615]+y[615]+z[615]);
assign {c[617],s[616]} = (x[616]+y[616]+z[616]);
assign {c[618],s[617]} = (x[617]+y[617]+z[617]);
assign {c[619],s[618]} = (x[618]+y[618]+z[618]);
assign {c[620],s[619]} = (x[619]+y[619]+z[619]);
assign {c[621],s[620]} = (x[620]+y[620]+z[620]);
assign {c[622],s[621]} = (x[621]+y[621]+z[621]);
assign {c[623],s[622]} = (x[622]+y[622]+z[622]);
assign {c[624],s[623]} = (x[623]+y[623]+z[623]);
assign {c[625],s[624]} = (x[624]+y[624]+z[624]);
assign {c[626],s[625]} = (x[625]+y[625]+z[625]);
assign {c[627],s[626]} = (x[626]+y[626]+z[626]);
assign {c[628],s[627]} = (x[627]+y[627]+z[627]);
assign {c[629],s[628]} = (x[628]+y[628]+z[628]);
assign {c[630],s[629]} = (x[629]+y[629]+z[629]);
assign {c[631],s[630]} = (x[630]+y[630]+z[630]);
assign {c[632],s[631]} = (x[631]+y[631]+z[631]);
assign {c[633],s[632]} = (x[632]+y[632]+z[632]);
assign {c[634],s[633]} = (x[633]+y[633]+z[633]);
assign {c[635],s[634]} = (x[634]+y[634]+z[634]);
assign {c[636],s[635]} = (x[635]+y[635]+z[635]);
assign {c[637],s[636]} = (x[636]+y[636]+z[636]);
assign {c[638],s[637]} = (x[637]+y[637]+z[637]);
assign {c[639],s[638]} = (x[638]+y[638]+z[638]);
assign {c[640],s[639]} = (x[639]+y[639]+z[639]);
assign {c[641],s[640]} = (x[640]+y[640]+z[640]);
assign {c[642],s[641]} = (x[641]+y[641]+z[641]);
assign {c[643],s[642]} = (x[642]+y[642]+z[642]);
assign {c[644],s[643]} = (x[643]+y[643]+z[643]);
assign {c[645],s[644]} = (x[644]+y[644]+z[644]);
assign {c[646],s[645]} = (x[645]+y[645]+z[645]);
assign {c[647],s[646]} = (x[646]+y[646]+z[646]);
assign {c[648],s[647]} = (x[647]+y[647]+z[647]);
assign {c[649],s[648]} = (x[648]+y[648]+z[648]);
assign {c[650],s[649]} = (x[649]+y[649]+z[649]);
assign {c[651],s[650]} = (x[650]+y[650]+z[650]);
assign {c[652],s[651]} = (x[651]+y[651]+z[651]);
assign {c[653],s[652]} = (x[652]+y[652]+z[652]);
assign {c[654],s[653]} = (x[653]+y[653]+z[653]);
assign {c[655],s[654]} = (x[654]+y[654]+z[654]);
assign {c[656],s[655]} = (x[655]+y[655]+z[655]);
assign {c[657],s[656]} = (x[656]+y[656]+z[656]);
assign {c[658],s[657]} = (x[657]+y[657]+z[657]);
assign {c[659],s[658]} = (x[658]+y[658]+z[658]);
assign {c[660],s[659]} = (x[659]+y[659]+z[659]);
assign {c[661],s[660]} = (x[660]+y[660]+z[660]);
assign {c[662],s[661]} = (x[661]+y[661]+z[661]);
assign {c[663],s[662]} = (x[662]+y[662]+z[662]);
assign {c[664],s[663]} = (x[663]+y[663]+z[663]);
assign {c[665],s[664]} = (x[664]+y[664]+z[664]);
assign {c[666],s[665]} = (x[665]+y[665]+z[665]);
assign {c[667],s[666]} = (x[666]+y[666]+z[666]);
assign {c[668],s[667]} = (x[667]+y[667]+z[667]);
assign {c[669],s[668]} = (x[668]+y[668]+z[668]);
assign {c[670],s[669]} = (x[669]+y[669]+z[669]);
assign {c[671],s[670]} = (x[670]+y[670]+z[670]);
assign {c[672],s[671]} = (x[671]+y[671]+z[671]);
assign {c[673],s[672]} = (x[672]+y[672]+z[672]);
assign {c[674],s[673]} = (x[673]+y[673]+z[673]);
assign {c[675],s[674]} = (x[674]+y[674]+z[674]);
assign {c[676],s[675]} = (x[675]+y[675]+z[675]);
assign {c[677],s[676]} = (x[676]+y[676]+z[676]);
assign {c[678],s[677]} = (x[677]+y[677]+z[677]);
assign {c[679],s[678]} = (x[678]+y[678]+z[678]);
assign {c[680],s[679]} = (x[679]+y[679]+z[679]);
assign {c[681],s[680]} = (x[680]+y[680]+z[680]);
assign {c[682],s[681]} = (x[681]+y[681]+z[681]);
assign {c[683],s[682]} = (x[682]+y[682]+z[682]);
assign {c[684],s[683]} = (x[683]+y[683]+z[683]);
assign {c[685],s[684]} = (x[684]+y[684]+z[684]);
assign {c[686],s[685]} = (x[685]+y[685]+z[685]);
assign {c[687],s[686]} = (x[686]+y[686]+z[686]);
assign {c[688],s[687]} = (x[687]+y[687]+z[687]);
assign {c[689],s[688]} = (x[688]+y[688]+z[688]);
assign {c[690],s[689]} = (x[689]+y[689]+z[689]);
assign {c[691],s[690]} = (x[690]+y[690]+z[690]);
assign {c[692],s[691]} = (x[691]+y[691]+z[691]);
assign {c[693],s[692]} = (x[692]+y[692]+z[692]);
assign {c[694],s[693]} = (x[693]+y[693]+z[693]);
assign {c[695],s[694]} = (x[694]+y[694]+z[694]);
assign {c[696],s[695]} = (x[695]+y[695]+z[695]);
assign {c[697],s[696]} = (x[696]+y[696]+z[696]);
assign {c[698],s[697]} = (x[697]+y[697]+z[697]);
assign {c[699],s[698]} = (x[698]+y[698]+z[698]);
assign {c[700],s[699]} = (x[699]+y[699]+z[699]);
assign {c[701],s[700]} = (x[700]+y[700]+z[700]);
assign {c[702],s[701]} = (x[701]+y[701]+z[701]);
assign {c[703],s[702]} = (x[702]+y[702]+z[702]);
assign {c[704],s[703]} = (x[703]+y[703]+z[703]);
assign {c[705],s[704]} = (x[704]+y[704]+z[704]);
assign {c[706],s[705]} = (x[705]+y[705]+z[705]);
assign {c[707],s[706]} = (x[706]+y[706]+z[706]);
assign {c[708],s[707]} = (x[707]+y[707]+z[707]);
assign {c[709],s[708]} = (x[708]+y[708]+z[708]);
assign {c[710],s[709]} = (x[709]+y[709]+z[709]);
assign {c[711],s[710]} = (x[710]+y[710]+z[710]);
assign {c[712],s[711]} = (x[711]+y[711]+z[711]);
assign {c[713],s[712]} = (x[712]+y[712]+z[712]);
assign {c[714],s[713]} = (x[713]+y[713]+z[713]);
assign {c[715],s[714]} = (x[714]+y[714]+z[714]);
assign {c[716],s[715]} = (x[715]+y[715]+z[715]);
assign {c[717],s[716]} = (x[716]+y[716]+z[716]);
assign {c[718],s[717]} = (x[717]+y[717]+z[717]);
assign {c[719],s[718]} = (x[718]+y[718]+z[718]);
assign {c[720],s[719]} = (x[719]+y[719]+z[719]);
assign {c[721],s[720]} = (x[720]+y[720]+z[720]);
assign {c[722],s[721]} = (x[721]+y[721]+z[721]);
assign {c[723],s[722]} = (x[722]+y[722]+z[722]);
assign {c[724],s[723]} = (x[723]+y[723]+z[723]);
assign {c[725],s[724]} = (x[724]+y[724]+z[724]);
assign {c[726],s[725]} = (x[725]+y[725]+z[725]);
assign {c[727],s[726]} = (x[726]+y[726]+z[726]);
assign {c[728],s[727]} = (x[727]+y[727]+z[727]);
assign {c[729],s[728]} = (x[728]+y[728]+z[728]);
assign {c[730],s[729]} = (x[729]+y[729]+z[729]);
assign {c[731],s[730]} = (x[730]+y[730]+z[730]);
assign {c[732],s[731]} = (x[731]+y[731]+z[731]);
assign {c[733],s[732]} = (x[732]+y[732]+z[732]);
assign {c[734],s[733]} = (x[733]+y[733]+z[733]);
assign {c[735],s[734]} = (x[734]+y[734]+z[734]);
assign {c[736],s[735]} = (x[735]+y[735]+z[735]);
assign {c[737],s[736]} = (x[736]+y[736]+z[736]);
assign {c[738],s[737]} = (x[737]+y[737]+z[737]);
assign {c[739],s[738]} = (x[738]+y[738]+z[738]);
assign {c[740],s[739]} = (x[739]+y[739]+z[739]);
assign {c[741],s[740]} = (x[740]+y[740]+z[740]);
assign {c[742],s[741]} = (x[741]+y[741]+z[741]);
assign {c[743],s[742]} = (x[742]+y[742]+z[742]);
assign {c[744],s[743]} = (x[743]+y[743]+z[743]);
assign {c[745],s[744]} = (x[744]+y[744]+z[744]);
assign {c[746],s[745]} = (x[745]+y[745]+z[745]);
assign {c[747],s[746]} = (x[746]+y[746]+z[746]);
assign {c[748],s[747]} = (x[747]+y[747]+z[747]);
assign {c[749],s[748]} = (x[748]+y[748]+z[748]);
assign {c[750],s[749]} = (x[749]+y[749]+z[749]);
assign {c[751],s[750]} = (x[750]+y[750]+z[750]);
assign {c[752],s[751]} = (x[751]+y[751]+z[751]);
assign {c[753],s[752]} = (x[752]+y[752]+z[752]);
assign {c[754],s[753]} = (x[753]+y[753]+z[753]);
assign {c[755],s[754]} = (x[754]+y[754]+z[754]);
assign {c[756],s[755]} = (x[755]+y[755]+z[755]);
assign {c[757],s[756]} = (x[756]+y[756]+z[756]);
assign {c[758],s[757]} = (x[757]+y[757]+z[757]);
assign {c[759],s[758]} = (x[758]+y[758]+z[758]);
assign {c[760],s[759]} = (x[759]+y[759]+z[759]);
assign {c[761],s[760]} = (x[760]+y[760]+z[760]);
assign {c[762],s[761]} = (x[761]+y[761]+z[761]);
assign {c[763],s[762]} = (x[762]+y[762]+z[762]);
assign {c[764],s[763]} = (x[763]+y[763]+z[763]);
assign {c[765],s[764]} = (x[764]+y[764]+z[764]);
assign {c[766],s[765]} = (x[765]+y[765]+z[765]);
assign {c[767],s[766]} = (x[766]+y[766]+z[766]);
assign {c[768],s[767]} = (x[767]+y[767]+z[767]);
assign {c[769],s[768]} = (x[768]+y[768]+z[768]);
assign {c[770],s[769]} = (x[769]+y[769]+z[769]);
assign {c[771],s[770]} = (x[770]+y[770]+z[770]);
assign {c[772],s[771]} = (x[771]+y[771]+z[771]);
assign {c[773],s[772]} = (x[772]+y[772]+z[772]);
assign {c[774],s[773]} = (x[773]+y[773]+z[773]);
assign {c[775],s[774]} = (x[774]+y[774]+z[774]);
assign {c[776],s[775]} = (x[775]+y[775]+z[775]);
assign {c[777],s[776]} = (x[776]+y[776]+z[776]);
assign {c[778],s[777]} = (x[777]+y[777]+z[777]);
assign {c[779],s[778]} = (x[778]+y[778]+z[778]);
assign {c[780],s[779]} = (x[779]+y[779]+z[779]);
assign {c[781],s[780]} = (x[780]+y[780]+z[780]);
assign {c[782],s[781]} = (x[781]+y[781]+z[781]);
assign {c[783],s[782]} = (x[782]+y[782]+z[782]);
assign {c[784],s[783]} = (x[783]+y[783]+z[783]);
assign {c[785],s[784]} = (x[784]+y[784]+z[784]);
assign {c[786],s[785]} = (x[785]+y[785]+z[785]);
assign {c[787],s[786]} = (x[786]+y[786]+z[786]);
assign {c[788],s[787]} = (x[787]+y[787]+z[787]);
assign {c[789],s[788]} = (x[788]+y[788]+z[788]);
assign {c[790],s[789]} = (x[789]+y[789]+z[789]);
assign {c[791],s[790]} = (x[790]+y[790]+z[790]);
assign {c[792],s[791]} = (x[791]+y[791]+z[791]);
assign {c[793],s[792]} = (x[792]+y[792]+z[792]);
assign {c[794],s[793]} = (x[793]+y[793]+z[793]);
assign {c[795],s[794]} = (x[794]+y[794]+z[794]);
assign {c[796],s[795]} = (x[795]+y[795]+z[795]);
assign {c[797],s[796]} = (x[796]+y[796]+z[796]);
assign {c[798],s[797]} = (x[797]+y[797]+z[797]);
assign {c[799],s[798]} = (x[798]+y[798]+z[798]);
assign {c[800],s[799]} = (x[799]+y[799]+z[799]);
assign {c[801],s[800]} = (x[800]+y[800]+z[800]);
assign {c[802],s[801]} = (x[801]+y[801]+z[801]);
assign {c[803],s[802]} = (x[802]+y[802]+z[802]);
assign {c[804],s[803]} = (x[803]+y[803]+z[803]);
assign {c[805],s[804]} = (x[804]+y[804]+z[804]);
assign {c[806],s[805]} = (x[805]+y[805]+z[805]);
assign {c[807],s[806]} = (x[806]+y[806]+z[806]);
assign {c[808],s[807]} = (x[807]+y[807]+z[807]);
assign {c[809],s[808]} = (x[808]+y[808]+z[808]);
assign {c[810],s[809]} = (x[809]+y[809]+z[809]);
assign {c[811],s[810]} = (x[810]+y[810]+z[810]);
assign {c[812],s[811]} = (x[811]+y[811]+z[811]);
assign {c[813],s[812]} = (x[812]+y[812]+z[812]);
assign {c[814],s[813]} = (x[813]+y[813]+z[813]);
assign {c[815],s[814]} = (x[814]+y[814]+z[814]);
assign {c[816],s[815]} = (x[815]+y[815]+z[815]);
assign {c[817],s[816]} = (x[816]+y[816]+z[816]);
assign {c[818],s[817]} = (x[817]+y[817]+z[817]);
assign {c[819],s[818]} = (x[818]+y[818]+z[818]);
assign {c[820],s[819]} = (x[819]+y[819]+z[819]);
assign {c[821],s[820]} = (x[820]+y[820]+z[820]);
assign {c[822],s[821]} = (x[821]+y[821]+z[821]);
assign {c[823],s[822]} = (x[822]+y[822]+z[822]);
assign {c[824],s[823]} = (x[823]+y[823]+z[823]);
assign {c[825],s[824]} = (x[824]+y[824]+z[824]);
assign {c[826],s[825]} = (x[825]+y[825]+z[825]);
assign {c[827],s[826]} = (x[826]+y[826]+z[826]);
assign {c[828],s[827]} = (x[827]+y[827]+z[827]);
assign {c[829],s[828]} = (x[828]+y[828]+z[828]);
assign {c[830],s[829]} = (x[829]+y[829]+z[829]);
assign {c[831],s[830]} = (x[830]+y[830]+z[830]);
assign {c[832],s[831]} = (x[831]+y[831]+z[831]);
assign {c[833],s[832]} = (x[832]+y[832]+z[832]);
assign {c[834],s[833]} = (x[833]+y[833]+z[833]);
assign {c[835],s[834]} = (x[834]+y[834]+z[834]);
assign {c[836],s[835]} = (x[835]+y[835]+z[835]);
assign {c[837],s[836]} = (x[836]+y[836]+z[836]);
assign {c[838],s[837]} = (x[837]+y[837]+z[837]);
assign {c[839],s[838]} = (x[838]+y[838]+z[838]);
assign {c[840],s[839]} = (x[839]+y[839]+z[839]);
assign {c[841],s[840]} = (x[840]+y[840]+z[840]);
assign {c[842],s[841]} = (x[841]+y[841]+z[841]);
assign {c[843],s[842]} = (x[842]+y[842]+z[842]);
assign {c[844],s[843]} = (x[843]+y[843]+z[843]);
assign {c[845],s[844]} = (x[844]+y[844]+z[844]);
assign {c[846],s[845]} = (x[845]+y[845]+z[845]);
assign {c[847],s[846]} = (x[846]+y[846]+z[846]);
assign {c[848],s[847]} = (x[847]+y[847]+z[847]);
assign {c[849],s[848]} = (x[848]+y[848]+z[848]);
assign {c[850],s[849]} = (x[849]+y[849]+z[849]);
assign {c[851],s[850]} = (x[850]+y[850]+z[850]);
assign {c[852],s[851]} = (x[851]+y[851]+z[851]);
assign {c[853],s[852]} = (x[852]+y[852]+z[852]);
assign {c[854],s[853]} = (x[853]+y[853]+z[853]);
assign {c[855],s[854]} = (x[854]+y[854]+z[854]);
assign {c[856],s[855]} = (x[855]+y[855]+z[855]);
assign {c[857],s[856]} = (x[856]+y[856]+z[856]);
assign {c[858],s[857]} = (x[857]+y[857]+z[857]);
assign {c[859],s[858]} = (x[858]+y[858]+z[858]);
assign {c[860],s[859]} = (x[859]+y[859]+z[859]);
assign {c[861],s[860]} = (x[860]+y[860]+z[860]);
assign {c[862],s[861]} = (x[861]+y[861]+z[861]);
assign {c[863],s[862]} = (x[862]+y[862]+z[862]);
assign {c[864],s[863]} = (x[863]+y[863]+z[863]);
assign {c[865],s[864]} = (x[864]+y[864]+z[864]);
assign {c[866],s[865]} = (x[865]+y[865]+z[865]);
assign {c[867],s[866]} = (x[866]+y[866]+z[866]);
assign {c[868],s[867]} = (x[867]+y[867]+z[867]);
assign {c[869],s[868]} = (x[868]+y[868]+z[868]);
assign {c[870],s[869]} = (x[869]+y[869]+z[869]);
assign {c[871],s[870]} = (x[870]+y[870]+z[870]);
assign {c[872],s[871]} = (x[871]+y[871]+z[871]);
assign {c[873],s[872]} = (x[872]+y[872]+z[872]);
assign {c[874],s[873]} = (x[873]+y[873]+z[873]);
assign {c[875],s[874]} = (x[874]+y[874]+z[874]);
assign {c[876],s[875]} = (x[875]+y[875]+z[875]);
assign {c[877],s[876]} = (x[876]+y[876]+z[876]);
assign {c[878],s[877]} = (x[877]+y[877]+z[877]);
assign {c[879],s[878]} = (x[878]+y[878]+z[878]);
assign {c[880],s[879]} = (x[879]+y[879]+z[879]);
assign {c[881],s[880]} = (x[880]+y[880]+z[880]);
assign {c[882],s[881]} = (x[881]+y[881]+z[881]);
assign {c[883],s[882]} = (x[882]+y[882]+z[882]);
assign {c[884],s[883]} = (x[883]+y[883]+z[883]);
assign {c[885],s[884]} = (x[884]+y[884]+z[884]);
assign {c[886],s[885]} = (x[885]+y[885]+z[885]);
assign {c[887],s[886]} = (x[886]+y[886]+z[886]);
assign {c[888],s[887]} = (x[887]+y[887]+z[887]);
assign {c[889],s[888]} = (x[888]+y[888]+z[888]);
assign {c[890],s[889]} = (x[889]+y[889]+z[889]);
assign {c[891],s[890]} = (x[890]+y[890]+z[890]);
assign {c[892],s[891]} = (x[891]+y[891]+z[891]);
assign {c[893],s[892]} = (x[892]+y[892]+z[892]);
assign {c[894],s[893]} = (x[893]+y[893]+z[893]);
assign {c[895],s[894]} = (x[894]+y[894]+z[894]);
assign {c[896],s[895]} = (x[895]+y[895]+z[895]);
assign {c[897],s[896]} = (x[896]+y[896]+z[896]);
assign {c[898],s[897]} = (x[897]+y[897]+z[897]);
assign {c[899],s[898]} = (x[898]+y[898]+z[898]);
assign {c[900],s[899]} = (x[899]+y[899]+z[899]);
assign {c[901],s[900]} = (x[900]+y[900]+z[900]);
assign {c[902],s[901]} = (x[901]+y[901]+z[901]);
assign {c[903],s[902]} = (x[902]+y[902]+z[902]);
assign {c[904],s[903]} = (x[903]+y[903]+z[903]);
assign {c[905],s[904]} = (x[904]+y[904]+z[904]);
assign {c[906],s[905]} = (x[905]+y[905]+z[905]);
assign {c[907],s[906]} = (x[906]+y[906]+z[906]);
assign {c[908],s[907]} = (x[907]+y[907]+z[907]);
assign {c[909],s[908]} = (x[908]+y[908]+z[908]);
assign {c[910],s[909]} = (x[909]+y[909]+z[909]);
assign {c[911],s[910]} = (x[910]+y[910]+z[910]);
assign {c[912],s[911]} = (x[911]+y[911]+z[911]);
assign {c[913],s[912]} = (x[912]+y[912]+z[912]);
assign {c[914],s[913]} = (x[913]+y[913]+z[913]);
assign {c[915],s[914]} = (x[914]+y[914]+z[914]);
assign {c[916],s[915]} = (x[915]+y[915]+z[915]);
assign {c[917],s[916]} = (x[916]+y[916]+z[916]);
assign {c[918],s[917]} = (x[917]+y[917]+z[917]);
assign {c[919],s[918]} = (x[918]+y[918]+z[918]);
assign {c[920],s[919]} = (x[919]+y[919]+z[919]);
assign {c[921],s[920]} = (x[920]+y[920]+z[920]);
assign {c[922],s[921]} = (x[921]+y[921]+z[921]);
assign {c[923],s[922]} = (x[922]+y[922]+z[922]);
assign {c[924],s[923]} = (x[923]+y[923]+z[923]);
assign {c[925],s[924]} = (x[924]+y[924]+z[924]);
assign {c[926],s[925]} = (x[925]+y[925]+z[925]);
assign {c[927],s[926]} = (x[926]+y[926]+z[926]);
assign {c[928],s[927]} = (x[927]+y[927]+z[927]);
assign {c[929],s[928]} = (x[928]+y[928]+z[928]);
assign {c[930],s[929]} = (x[929]+y[929]+z[929]);
assign {c[931],s[930]} = (x[930]+y[930]+z[930]);
assign {c[932],s[931]} = (x[931]+y[931]+z[931]);
assign {c[933],s[932]} = (x[932]+y[932]+z[932]);
assign {c[934],s[933]} = (x[933]+y[933]+z[933]);
assign {c[935],s[934]} = (x[934]+y[934]+z[934]);
assign {c[936],s[935]} = (x[935]+y[935]+z[935]);
assign {c[937],s[936]} = (x[936]+y[936]+z[936]);
assign {c[938],s[937]} = (x[937]+y[937]+z[937]);
assign {c[939],s[938]} = (x[938]+y[938]+z[938]);
assign {c[940],s[939]} = (x[939]+y[939]+z[939]);
assign {c[941],s[940]} = (x[940]+y[940]+z[940]);
assign {c[942],s[941]} = (x[941]+y[941]+z[941]);
assign {c[943],s[942]} = (x[942]+y[942]+z[942]);
assign {c[944],s[943]} = (x[943]+y[943]+z[943]);
assign {c[945],s[944]} = (x[944]+y[944]+z[944]);
assign {c[946],s[945]} = (x[945]+y[945]+z[945]);
assign {c[947],s[946]} = (x[946]+y[946]+z[946]);
assign {c[948],s[947]} = (x[947]+y[947]+z[947]);
assign {c[949],s[948]} = (x[948]+y[948]+z[948]);
assign {c[950],s[949]} = (x[949]+y[949]+z[949]);
assign {c[951],s[950]} = (x[950]+y[950]+z[950]);
assign {c[952],s[951]} = (x[951]+y[951]+z[951]);
assign {c[953],s[952]} = (x[952]+y[952]+z[952]);
assign {c[954],s[953]} = (x[953]+y[953]+z[953]);
assign {c[955],s[954]} = (x[954]+y[954]+z[954]);
assign {c[956],s[955]} = (x[955]+y[955]+z[955]);
assign {c[957],s[956]} = (x[956]+y[956]+z[956]);
assign {c[958],s[957]} = (x[957]+y[957]+z[957]);
assign {c[959],s[958]} = (x[958]+y[958]+z[958]);
assign {c[960],s[959]} = (x[959]+y[959]+z[959]);
assign {c[961],s[960]} = (x[960]+y[960]+z[960]);
assign {c[962],s[961]} = (x[961]+y[961]+z[961]);
assign {c[963],s[962]} = (x[962]+y[962]+z[962]);
assign {c[964],s[963]} = (x[963]+y[963]+z[963]);
assign {c[965],s[964]} = (x[964]+y[964]+z[964]);
assign {c[966],s[965]} = (x[965]+y[965]+z[965]);
assign {c[967],s[966]} = (x[966]+y[966]+z[966]);
assign {c[968],s[967]} = (x[967]+y[967]+z[967]);
assign {c[969],s[968]} = (x[968]+y[968]+z[968]);
assign {c[970],s[969]} = (x[969]+y[969]+z[969]);
assign {c[971],s[970]} = (x[970]+y[970]+z[970]);
assign {c[972],s[971]} = (x[971]+y[971]+z[971]);
assign {c[973],s[972]} = (x[972]+y[972]+z[972]);
assign {c[974],s[973]} = (x[973]+y[973]+z[973]);
assign {c[975],s[974]} = (x[974]+y[974]+z[974]);
assign {c[976],s[975]} = (x[975]+y[975]+z[975]);
assign {c[977],s[976]} = (x[976]+y[976]+z[976]);
assign {c[978],s[977]} = (x[977]+y[977]+z[977]);
assign {c[979],s[978]} = (x[978]+y[978]+z[978]);
assign {c[980],s[979]} = (x[979]+y[979]+z[979]);
assign {c[981],s[980]} = (x[980]+y[980]+z[980]);
assign {c[982],s[981]} = (x[981]+y[981]+z[981]);
assign {c[983],s[982]} = (x[982]+y[982]+z[982]);
assign {c[984],s[983]} = (x[983]+y[983]+z[983]);
assign {c[985],s[984]} = (x[984]+y[984]+z[984]);
assign {c[986],s[985]} = (x[985]+y[985]+z[985]);
assign {c[987],s[986]} = (x[986]+y[986]+z[986]);
assign {c[988],s[987]} = (x[987]+y[987]+z[987]);
assign {c[989],s[988]} = (x[988]+y[988]+z[988]);
assign {c[990],s[989]} = (x[989]+y[989]+z[989]);
assign {c[991],s[990]} = (x[990]+y[990]+z[990]);
assign {c[992],s[991]} = (x[991]+y[991]+z[991]);
assign {c[993],s[992]} = (x[992]+y[992]+z[992]);
assign {c[994],s[993]} = (x[993]+y[993]+z[993]);
assign {c[995],s[994]} = (x[994]+y[994]+z[994]);
assign {c[996],s[995]} = (x[995]+y[995]+z[995]);
assign {c[997],s[996]} = (x[996]+y[996]+z[996]);
assign {c[998],s[997]} = (x[997]+y[997]+z[997]);
assign {c[999],s[998]} = (x[998]+y[998]+z[998]);
assign {c[1000],s[999]} = (x[999]+y[999]+z[999]);
assign {c[1001],s[1000]} = (x[1000]+y[1000]+z[1000]);
assign {c[1002],s[1001]} = (x[1001]+y[1001]+z[1001]);
assign {c[1003],s[1002]} = (x[1002]+y[1002]+z[1002]);
assign {c[1004],s[1003]} = (x[1003]+y[1003]+z[1003]);
assign {c[1005],s[1004]} = (x[1004]+y[1004]+z[1004]);
assign {c[1006],s[1005]} = (x[1005]+y[1005]+z[1005]);
assign {c[1007],s[1006]} = (x[1006]+y[1006]+z[1006]);
assign {c[1008],s[1007]} = (x[1007]+y[1007]+z[1007]);
assign {c[1009],s[1008]} = (x[1008]+y[1008]+z[1008]);
assign {c[1010],s[1009]} = (x[1009]+y[1009]+z[1009]);
assign {c[1011],s[1010]} = (x[1010]+y[1010]+z[1010]);
assign {c[1012],s[1011]} = (x[1011]+y[1011]+z[1011]);
assign {c[1013],s[1012]} = (x[1012]+y[1012]+z[1012]);
assign {c[1014],s[1013]} = (x[1013]+y[1013]+z[1013]);
assign {c[1015],s[1014]} = (x[1014]+y[1014]+z[1014]);
assign {c[1016],s[1015]} = (x[1015]+y[1015]+z[1015]);
assign {c[1017],s[1016]} = (x[1016]+y[1016]+z[1016]);
assign {c[1018],s[1017]} = (x[1017]+y[1017]+z[1017]);
assign {c[1019],s[1018]} = (x[1018]+y[1018]+z[1018]);
assign {c[1020],s[1019]} = (x[1019]+y[1019]+z[1019]);
assign {c[1021],s[1020]} = (x[1020]+y[1020]+z[1020]);
assign {c[1022],s[1021]} = (x[1021]+y[1021]+z[1021]);
assign {c[1023],s[1022]} = (x[1022]+y[1022]+z[1022]);
assign {c[1024],s[1023]} = (x[1023]+y[1023]+z[1023]);
assign {c[1025],s[1024]} = (x[1024]+y[1024]+z[1024]);
assign {c[1026],s[1025]} = (x[1025]+y[1025]+z[1025]);
assign {c[1027],s[1026]} = (x[1026]+y[1026]+z[1026]);
assign {c[1028],s[1027]} = (x[1027]+y[1027]+z[1027]);
assign {c[1029],s[1028]} = (x[1028]+y[1028]+z[1028]);
assign {c[1030],s[1029]} = (x[1029]+y[1029]+z[1029]);
assign {c[1031],s[1030]} = (x[1030]+y[1030]+z[1030]);
assign {c[1032],s[1031]} = (x[1031]+y[1031]+z[1031]);
assign {c[1033],s[1032]} = (x[1032]+y[1032]+z[1032]);
assign {c[1034],s[1033]} = (x[1033]+y[1033]+z[1033]);
assign {c[1035],s[1034]} = (x[1034]+y[1034]+z[1034]);
assign {c[1036],s[1035]} = (x[1035]+y[1035]+z[1035]);
assign {c[1037],s[1036]} = (x[1036]+y[1036]+z[1036]);
assign {c[1038],s[1037]} = (x[1037]+y[1037]+z[1037]);
assign {c[1039],s[1038]} = (x[1038]+y[1038]+z[1038]);
assign {c[1040],s[1039]} = (x[1039]+y[1039]+z[1039]);
assign {c[1041],s[1040]} = (x[1040]+y[1040]+z[1040]);
assign {c[1042],s[1041]} = (x[1041]+y[1041]+z[1041]);
assign {c[1043],s[1042]} = (x[1042]+y[1042]+z[1042]);
assign {c[1044],s[1043]} = (x[1043]+y[1043]+z[1043]);
assign {c[1045],s[1044]} = (x[1044]+y[1044]+z[1044]);
assign {c[1046],s[1045]} = (x[1045]+y[1045]+z[1045]);
assign {c[1047],s[1046]} = (x[1046]+y[1046]+z[1046]);
assign {c[1048],s[1047]} = (x[1047]+y[1047]+z[1047]);
assign {c[1049],s[1048]} = (x[1048]+y[1048]+z[1048]);
assign {c[1050],s[1049]} = (x[1049]+y[1049]+z[1049]);
assign {c[1051],s[1050]} = (x[1050]+y[1050]+z[1050]);
assign {c[1052],s[1051]} = (x[1051]+y[1051]+z[1051]);
assign {c[1053],s[1052]} = (x[1052]+y[1052]+z[1052]);
assign {c[1054],s[1053]} = (x[1053]+y[1053]+z[1053]);
assign {c[1055],s[1054]} = (x[1054]+y[1054]+z[1054]);
assign {c[1056],s[1055]} = (x[1055]+y[1055]+z[1055]);
assign {c[1057],s[1056]} = (x[1056]+y[1056]+z[1056]);
assign {c[1058],s[1057]} = (x[1057]+y[1057]+z[1057]);
assign {c[1059],s[1058]} = (x[1058]+y[1058]+z[1058]);
assign {c[1060],s[1059]} = (x[1059]+y[1059]+z[1059]);
assign {c[1061],s[1060]} = (x[1060]+y[1060]+z[1060]);
assign {c[1062],s[1061]} = (x[1061]+y[1061]+z[1061]);
assign {c[1063],s[1062]} = (x[1062]+y[1062]+z[1062]);
assign {c[1064],s[1063]} = (x[1063]+y[1063]+z[1063]);
assign {c[1065],s[1064]} = (x[1064]+y[1064]+z[1064]);
assign {c[1066],s[1065]} = (x[1065]+y[1065]+z[1065]);
assign {c[1067],s[1066]} = (x[1066]+y[1066]+z[1066]);
assign {c[1068],s[1067]} = (x[1067]+y[1067]+z[1067]);
assign {c[1069],s[1068]} = (x[1068]+y[1068]+z[1068]);
assign {c[1070],s[1069]} = (x[1069]+y[1069]+z[1069]);
assign {c[1071],s[1070]} = (x[1070]+y[1070]+z[1070]);
assign {c[1072],s[1071]} = (x[1071]+y[1071]+z[1071]);
assign {c[1073],s[1072]} = (x[1072]+y[1072]+z[1072]);
assign {c[1074],s[1073]} = (x[1073]+y[1073]+z[1073]);
assign {c[1075],s[1074]} = (x[1074]+y[1074]+z[1074]);
assign {c[1076],s[1075]} = (x[1075]+y[1075]+z[1075]);
assign {c[1077],s[1076]} = (x[1076]+y[1076]+z[1076]);
assign {c[1078],s[1077]} = (x[1077]+y[1077]+z[1077]);
assign {c[1079],s[1078]} = (x[1078]+y[1078]+z[1078]);
assign {c[1080],s[1079]} = (x[1079]+y[1079]+z[1079]);
assign {c[1081],s[1080]} = (x[1080]+y[1080]+z[1080]);
assign {c[1082],s[1081]} = (x[1081]+y[1081]+z[1081]);
assign {c[1083],s[1082]} = (x[1082]+y[1082]+z[1082]);
assign {c[1084],s[1083]} = (x[1083]+y[1083]+z[1083]);
assign {c[1085],s[1084]} = (x[1084]+y[1084]+z[1084]);
assign {c[1086],s[1085]} = (x[1085]+y[1085]+z[1085]);
assign {c[1087],s[1086]} = (x[1086]+y[1086]+z[1086]);
assign {c[1088],s[1087]} = (x[1087]+y[1087]+z[1087]);
assign {c[1089],s[1088]} = (x[1088]+y[1088]+z[1088]);
assign {c[1090],s[1089]} = (x[1089]+y[1089]+z[1089]);
assign {c[1091],s[1090]} = (x[1090]+y[1090]+z[1090]);
assign {c[1092],s[1091]} = (x[1091]+y[1091]+z[1091]);
assign {c[1093],s[1092]} = (x[1092]+y[1092]+z[1092]);
assign {c[1094],s[1093]} = (x[1093]+y[1093]+z[1093]);
assign {c[1095],s[1094]} = (x[1094]+y[1094]+z[1094]);
assign {c[1096],s[1095]} = (x[1095]+y[1095]+z[1095]);
assign {c[1097],s[1096]} = (x[1096]+y[1096]+z[1096]);
assign {c[1098],s[1097]} = (x[1097]+y[1097]+z[1097]);
assign {c[1099],s[1098]} = (x[1098]+y[1098]+z[1098]);
assign {c[1100],s[1099]} = (x[1099]+y[1099]+z[1099]);
assign {c[1101],s[1100]} = (x[1100]+y[1100]+z[1100]);
assign {c[1102],s[1101]} = (x[1101]+y[1101]+z[1101]);
assign {c[1103],s[1102]} = (x[1102]+y[1102]+z[1102]);
assign {c[1104],s[1103]} = (x[1103]+y[1103]+z[1103]);
assign {c[1105],s[1104]} = (x[1104]+y[1104]+z[1104]);
assign {c[1106],s[1105]} = (x[1105]+y[1105]+z[1105]);
assign {c[1107],s[1106]} = (x[1106]+y[1106]+z[1106]);
assign {c[1108],s[1107]} = (x[1107]+y[1107]+z[1107]);
assign {c[1109],s[1108]} = (x[1108]+y[1108]+z[1108]);
assign {c[1110],s[1109]} = (x[1109]+y[1109]+z[1109]);
assign {c[1111],s[1110]} = (x[1110]+y[1110]+z[1110]);
assign {c[1112],s[1111]} = (x[1111]+y[1111]+z[1111]);
assign {c[1113],s[1112]} = (x[1112]+y[1112]+z[1112]);
assign {c[1114],s[1113]} = (x[1113]+y[1113]+z[1113]);
assign {c[1115],s[1114]} = (x[1114]+y[1114]+z[1114]);
assign {c[1116],s[1115]} = (x[1115]+y[1115]+z[1115]);
assign {c[1117],s[1116]} = (x[1116]+y[1116]+z[1116]);
assign {c[1118],s[1117]} = (x[1117]+y[1117]+z[1117]);
assign {c[1119],s[1118]} = (x[1118]+y[1118]+z[1118]);
assign {c[1120],s[1119]} = (x[1119]+y[1119]+z[1119]);
assign {c[1121],s[1120]} = (x[1120]+y[1120]+z[1120]);
assign {c[1122],s[1121]} = (x[1121]+y[1121]+z[1121]);
assign {c[1123],s[1122]} = (x[1122]+y[1122]+z[1122]);
assign {c[1124],s[1123]} = (x[1123]+y[1123]+z[1123]);
assign {c[1125],s[1124]} = (x[1124]+y[1124]+z[1124]);
assign {c[1126],s[1125]} = (x[1125]+y[1125]+z[1125]);
assign {c[1127],s[1126]} = (x[1126]+y[1126]+z[1126]);
assign {c[1128],s[1127]} = (x[1127]+y[1127]+z[1127]);
assign {c[1129],s[1128]} = (x[1128]+y[1128]+z[1128]);
assign {c[1130],s[1129]} = (x[1129]+y[1129]+z[1129]);
assign {c[1131],s[1130]} = (x[1130]+y[1130]+z[1130]);
assign {c[1132],s[1131]} = (x[1131]+y[1131]+z[1131]);
assign {c[1133],s[1132]} = (x[1132]+y[1132]+z[1132]);
assign {c[1134],s[1133]} = (x[1133]+y[1133]+z[1133]);
assign {c[1135],s[1134]} = (x[1134]+y[1134]+z[1134]);
assign {c[1136],s[1135]} = (x[1135]+y[1135]+z[1135]);
assign {c[1137],s[1136]} = (x[1136]+y[1136]+z[1136]);
assign {c[1138],s[1137]} = (x[1137]+y[1137]+z[1137]);
assign {c[1139],s[1138]} = (x[1138]+y[1138]+z[1138]);
assign {c[1140],s[1139]} = (x[1139]+y[1139]+z[1139]);
assign {c[1141],s[1140]} = (x[1140]+y[1140]+z[1140]);
assign {c[1142],s[1141]} = (x[1141]+y[1141]+z[1141]);
assign {c[1143],s[1142]} = (x[1142]+y[1142]+z[1142]);
assign {c[1144],s[1143]} = (x[1143]+y[1143]+z[1143]);
assign {c[1145],s[1144]} = (x[1144]+y[1144]+z[1144]);
assign {c[1146],s[1145]} = (x[1145]+y[1145]+z[1145]);
assign {c[1147],s[1146]} = (x[1146]+y[1146]+z[1146]);
assign {c[1148],s[1147]} = (x[1147]+y[1147]+z[1147]);
assign {c[1149],s[1148]} = (x[1148]+y[1148]+z[1148]);
assign {c[1150],s[1149]} = (x[1149]+y[1149]+z[1149]);
assign {c[1151],s[1150]} = (x[1150]+y[1150]+z[1150]);
assign {c[1152],s[1151]} = (x[1151]+y[1151]+z[1151]);
assign {c[1153],s[1152]} = (x[1152]+y[1152]+z[1152]);
assign {c[1154],s[1153]} = (x[1153]+y[1153]+z[1153]);
assign {c[1155],s[1154]} = (x[1154]+y[1154]+z[1154]);
assign {c[1156],s[1155]} = (x[1155]+y[1155]+z[1155]);
assign {c[1157],s[1156]} = (x[1156]+y[1156]+z[1156]);
assign {c[1158],s[1157]} = (x[1157]+y[1157]+z[1157]);
assign {c[1159],s[1158]} = (x[1158]+y[1158]+z[1158]);
assign {c[1160],s[1159]} = (x[1159]+y[1159]+z[1159]);
assign {c[1161],s[1160]} = (x[1160]+y[1160]+z[1160]);
assign {c[1162],s[1161]} = (x[1161]+y[1161]+z[1161]);
assign {c[1163],s[1162]} = (x[1162]+y[1162]+z[1162]);
assign {c[1164],s[1163]} = (x[1163]+y[1163]+z[1163]);
assign {c[1165],s[1164]} = (x[1164]+y[1164]+z[1164]);
assign {c[1166],s[1165]} = (x[1165]+y[1165]+z[1165]);
assign {c[1167],s[1166]} = (x[1166]+y[1166]+z[1166]);
assign {c[1168],s[1167]} = (x[1167]+y[1167]+z[1167]);
assign {c[1169],s[1168]} = (x[1168]+y[1168]+z[1168]);
assign {c[1170],s[1169]} = (x[1169]+y[1169]+z[1169]);
assign {c[1171],s[1170]} = (x[1170]+y[1170]+z[1170]);
assign {c[1172],s[1171]} = (x[1171]+y[1171]+z[1171]);
assign {c[1173],s[1172]} = (x[1172]+y[1172]+z[1172]);
assign {c[1174],s[1173]} = (x[1173]+y[1173]+z[1173]);
assign {c[1175],s[1174]} = (x[1174]+y[1174]+z[1174]);
assign {c[1176],s[1175]} = (x[1175]+y[1175]+z[1175]);
assign {c[1177],s[1176]} = (x[1176]+y[1176]+z[1176]);
assign {c[1178],s[1177]} = (x[1177]+y[1177]+z[1177]);
assign {c[1179],s[1178]} = (x[1178]+y[1178]+z[1178]);
assign {c[1180],s[1179]} = (x[1179]+y[1179]+z[1179]);
assign {c[1181],s[1180]} = (x[1180]+y[1180]+z[1180]);
assign {c[1182],s[1181]} = (x[1181]+y[1181]+z[1181]);
assign {c[1183],s[1182]} = (x[1182]+y[1182]+z[1182]);
assign {c[1184],s[1183]} = (x[1183]+y[1183]+z[1183]);
assign {c[1185],s[1184]} = (x[1184]+y[1184]+z[1184]);
assign {c[1186],s[1185]} = (x[1185]+y[1185]+z[1185]);
assign {c[1187],s[1186]} = (x[1186]+y[1186]+z[1186]);
assign {c[1188],s[1187]} = (x[1187]+y[1187]+z[1187]);
assign {c[1189],s[1188]} = (x[1188]+y[1188]+z[1188]);
assign {c[1190],s[1189]} = (x[1189]+y[1189]+z[1189]);
assign {c[1191],s[1190]} = (x[1190]+y[1190]+z[1190]);
assign {c[1192],s[1191]} = (x[1191]+y[1191]+z[1191]);
assign {c[1193],s[1192]} = (x[1192]+y[1192]+z[1192]);
assign {c[1194],s[1193]} = (x[1193]+y[1193]+z[1193]);
assign {c[1195],s[1194]} = (x[1194]+y[1194]+z[1194]);
assign {c[1196],s[1195]} = (x[1195]+y[1195]+z[1195]);
assign {c[1197],s[1196]} = (x[1196]+y[1196]+z[1196]);
assign {c[1198],s[1197]} = (x[1197]+y[1197]+z[1197]);
assign {c[1199],s[1198]} = (x[1198]+y[1198]+z[1198]);
assign {c[1200],s[1199]} = (x[1199]+y[1199]+z[1199]);
assign {c[1201],s[1200]} = (x[1200]+y[1200]+z[1200]);
assign {c[1202],s[1201]} = (x[1201]+y[1201]+z[1201]);
assign {c[1203],s[1202]} = (x[1202]+y[1202]+z[1202]);
assign {c[1204],s[1203]} = (x[1203]+y[1203]+z[1203]);
assign {c[1205],s[1204]} = (x[1204]+y[1204]+z[1204]);
assign {c[1206],s[1205]} = (x[1205]+y[1205]+z[1205]);
assign {c[1207],s[1206]} = (x[1206]+y[1206]+z[1206]);
assign {c[1208],s[1207]} = (x[1207]+y[1207]+z[1207]);
assign {c[1209],s[1208]} = (x[1208]+y[1208]+z[1208]);
assign {c[1210],s[1209]} = (x[1209]+y[1209]+z[1209]);
assign {c[1211],s[1210]} = (x[1210]+y[1210]+z[1210]);
assign {c[1212],s[1211]} = (x[1211]+y[1211]+z[1211]);
assign {c[1213],s[1212]} = (x[1212]+y[1212]+z[1212]);
assign {c[1214],s[1213]} = (x[1213]+y[1213]+z[1213]);
assign {c[1215],s[1214]} = (x[1214]+y[1214]+z[1214]);
assign {c[1216],s[1215]} = (x[1215]+y[1215]+z[1215]);
assign {c[1217],s[1216]} = (x[1216]+y[1216]+z[1216]);
assign {c[1218],s[1217]} = (x[1217]+y[1217]+z[1217]);
assign {c[1219],s[1218]} = (x[1218]+y[1218]+z[1218]);
assign {c[1220],s[1219]} = (x[1219]+y[1219]+z[1219]);
assign {c[1221],s[1220]} = (x[1220]+y[1220]+z[1220]);
assign {c[1222],s[1221]} = (x[1221]+y[1221]+z[1221]);
assign {c[1223],s[1222]} = (x[1222]+y[1222]+z[1222]);
assign {c[1224],s[1223]} = (x[1223]+y[1223]+z[1223]);
assign {c[1225],s[1224]} = (x[1224]+y[1224]+z[1224]);
assign {c[1226],s[1225]} = (x[1225]+y[1225]+z[1225]);
assign {c[1227],s[1226]} = (x[1226]+y[1226]+z[1226]);
assign {c[1228],s[1227]} = (x[1227]+y[1227]+z[1227]);
assign {c[1229],s[1228]} = (x[1228]+y[1228]+z[1228]);
assign {c[1230],s[1229]} = (x[1229]+y[1229]+z[1229]);
assign {c[1231],s[1230]} = (x[1230]+y[1230]+z[1230]);
assign {c[1232],s[1231]} = (x[1231]+y[1231]+z[1231]);
assign {c[1233],s[1232]} = (x[1232]+y[1232]+z[1232]);
assign {c[1234],s[1233]} = (x[1233]+y[1233]+z[1233]);
assign {c[1235],s[1234]} = (x[1234]+y[1234]+z[1234]);
assign {c[1236],s[1235]} = (x[1235]+y[1235]+z[1235]);
assign {c[1237],s[1236]} = (x[1236]+y[1236]+z[1236]);
assign {c[1238],s[1237]} = (x[1237]+y[1237]+z[1237]);
assign {c[1239],s[1238]} = (x[1238]+y[1238]+z[1238]);
assign {c[1240],s[1239]} = (x[1239]+y[1239]+z[1239]);
assign {c[1241],s[1240]} = (x[1240]+y[1240]+z[1240]);
assign {c[1242],s[1241]} = (x[1241]+y[1241]+z[1241]);
assign {c[1243],s[1242]} = (x[1242]+y[1242]+z[1242]);
assign {c[1244],s[1243]} = (x[1243]+y[1243]+z[1243]);
assign {c[1245],s[1244]} = (x[1244]+y[1244]+z[1244]);
assign {c[1246],s[1245]} = (x[1245]+y[1245]+z[1245]);
assign {c[1247],s[1246]} = (x[1246]+y[1246]+z[1246]);
assign {c[1248],s[1247]} = (x[1247]+y[1247]+z[1247]);
assign {c[1249],s[1248]} = (x[1248]+y[1248]+z[1248]);
assign {c[1250],s[1249]} = (x[1249]+y[1249]+z[1249]);
assign {c[1251],s[1250]} = (x[1250]+y[1250]+z[1250]);
assign {c[1252],s[1251]} = (x[1251]+y[1251]+z[1251]);
assign {c[1253],s[1252]} = (x[1252]+y[1252]+z[1252]);
assign {c[1254],s[1253]} = (x[1253]+y[1253]+z[1253]);
assign {c[1255],s[1254]} = (x[1254]+y[1254]+z[1254]);
assign {c[1256],s[1255]} = (x[1255]+y[1255]+z[1255]);
assign {c[1257],s[1256]} = (x[1256]+y[1256]+z[1256]);
assign {c[1258],s[1257]} = (x[1257]+y[1257]+z[1257]);
assign {c[1259],s[1258]} = (x[1258]+y[1258]+z[1258]);
assign {c[1260],s[1259]} = (x[1259]+y[1259]+z[1259]);
assign {c[1261],s[1260]} = (x[1260]+y[1260]+z[1260]);
assign {c[1262],s[1261]} = (x[1261]+y[1261]+z[1261]);
assign {c[1263],s[1262]} = (x[1262]+y[1262]+z[1262]);
assign {c[1264],s[1263]} = (x[1263]+y[1263]+z[1263]);
assign {c[1265],s[1264]} = (x[1264]+y[1264]+z[1264]);
assign {c[1266],s[1265]} = (x[1265]+y[1265]+z[1265]);
assign {c[1267],s[1266]} = (x[1266]+y[1266]+z[1266]);
assign {c[1268],s[1267]} = (x[1267]+y[1267]+z[1267]);
assign {c[1269],s[1268]} = (x[1268]+y[1268]+z[1268]);
assign {c[1270],s[1269]} = (x[1269]+y[1269]+z[1269]);
assign {c[1271],s[1270]} = (x[1270]+y[1270]+z[1270]);
assign {c[1272],s[1271]} = (x[1271]+y[1271]+z[1271]);
assign {c[1273],s[1272]} = (x[1272]+y[1272]+z[1272]);
assign {c[1274],s[1273]} = (x[1273]+y[1273]+z[1273]);
assign {c[1275],s[1274]} = (x[1274]+y[1274]+z[1274]);
assign {c[1276],s[1275]} = (x[1275]+y[1275]+z[1275]);
assign {c[1277],s[1276]} = (x[1276]+y[1276]+z[1276]);
assign {c[1278],s[1277]} = (x[1277]+y[1277]+z[1277]);
assign {c[1279],s[1278]} = (x[1278]+y[1278]+z[1278]);
assign {c[1280],s[1279]} = (x[1279]+y[1279]+z[1279]);
assign {c[1281],s[1280]} = (x[1280]+y[1280]+z[1280]);
assign {c[1282],s[1281]} = (x[1281]+y[1281]+z[1281]);
assign {c[1283],s[1282]} = (x[1282]+y[1282]+z[1282]);
assign {c[1284],s[1283]} = (x[1283]+y[1283]+z[1283]);
assign {c[1285],s[1284]} = (x[1284]+y[1284]+z[1284]);
assign {c[1286],s[1285]} = (x[1285]+y[1285]+z[1285]);
assign {c[1287],s[1286]} = (x[1286]+y[1286]+z[1286]);
assign {c[1288],s[1287]} = (x[1287]+y[1287]+z[1287]);
assign {c[1289],s[1288]} = (x[1288]+y[1288]+z[1288]);
assign {c[1290],s[1289]} = (x[1289]+y[1289]+z[1289]);
assign {c[1291],s[1290]} = (x[1290]+y[1290]+z[1290]);
assign {c[1292],s[1291]} = (x[1291]+y[1291]+z[1291]);
assign {c[1293],s[1292]} = (x[1292]+y[1292]+z[1292]);
assign {c[1294],s[1293]} = (x[1293]+y[1293]+z[1293]);
assign {c[1295],s[1294]} = (x[1294]+y[1294]+z[1294]);
assign {c[1296],s[1295]} = (x[1295]+y[1295]+z[1295]);
assign {c[1297],s[1296]} = (x[1296]+y[1296]+z[1296]);
assign {c[1298],s[1297]} = (x[1297]+y[1297]+z[1297]);
assign {c[1299],s[1298]} = (x[1298]+y[1298]+z[1298]);
assign {c[1300],s[1299]} = (x[1299]+y[1299]+z[1299]);
assign {c[1301],s[1300]} = (x[1300]+y[1300]+z[1300]);
assign {c[1302],s[1301]} = (x[1301]+y[1301]+z[1301]);
assign {c[1303],s[1302]} = (x[1302]+y[1302]+z[1302]);
assign {c[1304],s[1303]} = (x[1303]+y[1303]+z[1303]);
assign {c[1305],s[1304]} = (x[1304]+y[1304]+z[1304]);
assign {c[1306],s[1305]} = (x[1305]+y[1305]+z[1305]);
assign {c[1307],s[1306]} = (x[1306]+y[1306]+z[1306]);
assign {c[1308],s[1307]} = (x[1307]+y[1307]+z[1307]);
assign {c[1309],s[1308]} = (x[1308]+y[1308]+z[1308]);
assign {c[1310],s[1309]} = (x[1309]+y[1309]+z[1309]);
assign {c[1311],s[1310]} = (x[1310]+y[1310]+z[1310]);
assign {c[1312],s[1311]} = (x[1311]+y[1311]+z[1311]);
assign {c[1313],s[1312]} = (x[1312]+y[1312]+z[1312]);
assign {c[1314],s[1313]} = (x[1313]+y[1313]+z[1313]);
assign {c[1315],s[1314]} = (x[1314]+y[1314]+z[1314]);
assign {c[1316],s[1315]} = (x[1315]+y[1315]+z[1315]);
assign {c[1317],s[1316]} = (x[1316]+y[1316]+z[1316]);
assign {c[1318],s[1317]} = (x[1317]+y[1317]+z[1317]);
assign {c[1319],s[1318]} = (x[1318]+y[1318]+z[1318]);
assign {c[1320],s[1319]} = (x[1319]+y[1319]+z[1319]);
assign {c[1321],s[1320]} = (x[1320]+y[1320]+z[1320]);
assign {c[1322],s[1321]} = (x[1321]+y[1321]+z[1321]);
assign {c[1323],s[1322]} = (x[1322]+y[1322]+z[1322]);
assign {c[1324],s[1323]} = (x[1323]+y[1323]+z[1323]);
assign {c[1325],s[1324]} = (x[1324]+y[1324]+z[1324]);
assign {c[1326],s[1325]} = (x[1325]+y[1325]+z[1325]);
assign {c[1327],s[1326]} = (x[1326]+y[1326]+z[1326]);
assign {c[1328],s[1327]} = (x[1327]+y[1327]+z[1327]);
assign {c[1329],s[1328]} = (x[1328]+y[1328]+z[1328]);
assign {c[1330],s[1329]} = (x[1329]+y[1329]+z[1329]);
assign {c[1331],s[1330]} = (x[1330]+y[1330]+z[1330]);
assign {c[1332],s[1331]} = (x[1331]+y[1331]+z[1331]);
assign {c[1333],s[1332]} = (x[1332]+y[1332]+z[1332]);
assign {c[1334],s[1333]} = (x[1333]+y[1333]+z[1333]);
assign {c[1335],s[1334]} = (x[1334]+y[1334]+z[1334]);
assign {c[1336],s[1335]} = (x[1335]+y[1335]+z[1335]);
assign {c[1337],s[1336]} = (x[1336]+y[1336]+z[1336]);
assign {c[1338],s[1337]} = (x[1337]+y[1337]+z[1337]);
assign {c[1339],s[1338]} = (x[1338]+y[1338]+z[1338]);
assign {c[1340],s[1339]} = (x[1339]+y[1339]+z[1339]);
assign {c[1341],s[1340]} = (x[1340]+y[1340]+z[1340]);
assign {c[1342],s[1341]} = (x[1341]+y[1341]+z[1341]);
assign {c[1343],s[1342]} = (x[1342]+y[1342]+z[1342]);
assign {c[1344],s[1343]} = (x[1343]+y[1343]+z[1343]);
assign {c[1345],s[1344]} = (x[1344]+y[1344]+z[1344]);
assign {c[1346],s[1345]} = (x[1345]+y[1345]+z[1345]);
assign {c[1347],s[1346]} = (x[1346]+y[1346]+z[1346]);
assign {c[1348],s[1347]} = (x[1347]+y[1347]+z[1347]);
assign {c[1349],s[1348]} = (x[1348]+y[1348]+z[1348]);
assign {c[1350],s[1349]} = (x[1349]+y[1349]+z[1349]);
assign {c[1351],s[1350]} = (x[1350]+y[1350]+z[1350]);
assign {c[1352],s[1351]} = (x[1351]+y[1351]+z[1351]);
assign {c[1353],s[1352]} = (x[1352]+y[1352]+z[1352]);
assign {c[1354],s[1353]} = (x[1353]+y[1353]+z[1353]);
assign {c[1355],s[1354]} = (x[1354]+y[1354]+z[1354]);
assign {c[1356],s[1355]} = (x[1355]+y[1355]+z[1355]);
assign {c[1357],s[1356]} = (x[1356]+y[1356]+z[1356]);
assign {c[1358],s[1357]} = (x[1357]+y[1357]+z[1357]);
assign {c[1359],s[1358]} = (x[1358]+y[1358]+z[1358]);
assign {c[1360],s[1359]} = (x[1359]+y[1359]+z[1359]);
assign {c[1361],s[1360]} = (x[1360]+y[1360]+z[1360]);
assign {c[1362],s[1361]} = (x[1361]+y[1361]+z[1361]);
assign {c[1363],s[1362]} = (x[1362]+y[1362]+z[1362]);
assign {c[1364],s[1363]} = (x[1363]+y[1363]+z[1363]);
assign {c[1365],s[1364]} = (x[1364]+y[1364]+z[1364]);
assign {c[1366],s[1365]} = (x[1365]+y[1365]+z[1365]);
assign {c[1367],s[1366]} = (x[1366]+y[1366]+z[1366]);
assign {c[1368],s[1367]} = (x[1367]+y[1367]+z[1367]);
assign {c[1369],s[1368]} = (x[1368]+y[1368]+z[1368]);
assign {c[1370],s[1369]} = (x[1369]+y[1369]+z[1369]);
assign {c[1371],s[1370]} = (x[1370]+y[1370]+z[1370]);
assign {c[1372],s[1371]} = (x[1371]+y[1371]+z[1371]);
assign {c[1373],s[1372]} = (x[1372]+y[1372]+z[1372]);
assign {c[1374],s[1373]} = (x[1373]+y[1373]+z[1373]);
assign {c[1375],s[1374]} = (x[1374]+y[1374]+z[1374]);
assign {c[1376],s[1375]} = (x[1375]+y[1375]+z[1375]);
assign {c[1377],s[1376]} = (x[1376]+y[1376]+z[1376]);
assign {c[1378],s[1377]} = (x[1377]+y[1377]+z[1377]);
assign {c[1379],s[1378]} = (x[1378]+y[1378]+z[1378]);
assign {c[1380],s[1379]} = (x[1379]+y[1379]+z[1379]);
assign {c[1381],s[1380]} = (x[1380]+y[1380]+z[1380]);
assign {c[1382],s[1381]} = (x[1381]+y[1381]+z[1381]);
assign {c[1383],s[1382]} = (x[1382]+y[1382]+z[1382]);
assign {c[1384],s[1383]} = (x[1383]+y[1383]+z[1383]);
assign {c[1385],s[1384]} = (x[1384]+y[1384]+z[1384]);
assign {c[1386],s[1385]} = (x[1385]+y[1385]+z[1385]);
assign {c[1387],s[1386]} = (x[1386]+y[1386]+z[1386]);
assign {c[1388],s[1387]} = (x[1387]+y[1387]+z[1387]);
assign {c[1389],s[1388]} = (x[1388]+y[1388]+z[1388]);
assign {c[1390],s[1389]} = (x[1389]+y[1389]+z[1389]);
assign {c[1391],s[1390]} = (x[1390]+y[1390]+z[1390]);
assign {c[1392],s[1391]} = (x[1391]+y[1391]+z[1391]);
assign {c[1393],s[1392]} = (x[1392]+y[1392]+z[1392]);
assign {c[1394],s[1393]} = (x[1393]+y[1393]+z[1393]);
assign {c[1395],s[1394]} = (x[1394]+y[1394]+z[1394]);
assign {c[1396],s[1395]} = (x[1395]+y[1395]+z[1395]);
assign {c[1397],s[1396]} = (x[1396]+y[1396]+z[1396]);
assign {c[1398],s[1397]} = (x[1397]+y[1397]+z[1397]);
assign {c[1399],s[1398]} = (x[1398]+y[1398]+z[1398]);
assign {c[1400],s[1399]} = (x[1399]+y[1399]+z[1399]);
assign {c[1401],s[1400]} = (x[1400]+y[1400]+z[1400]);
assign {c[1402],s[1401]} = (x[1401]+y[1401]+z[1401]);
assign {c[1403],s[1402]} = (x[1402]+y[1402]+z[1402]);
assign {c[1404],s[1403]} = (x[1403]+y[1403]+z[1403]);
assign {c[1405],s[1404]} = (x[1404]+y[1404]+z[1404]);
assign {c[1406],s[1405]} = (x[1405]+y[1405]+z[1405]);
assign {c[1407],s[1406]} = (x[1406]+y[1406]+z[1406]);
assign {c[1408],s[1407]} = (x[1407]+y[1407]+z[1407]);
assign {c[1409],s[1408]} = (x[1408]+y[1408]+z[1408]);
assign {c[1410],s[1409]} = (x[1409]+y[1409]+z[1409]);
assign {c[1411],s[1410]} = (x[1410]+y[1410]+z[1410]);
assign {c[1412],s[1411]} = (x[1411]+y[1411]+z[1411]);
assign {c[1413],s[1412]} = (x[1412]+y[1412]+z[1412]);
assign {c[1414],s[1413]} = (x[1413]+y[1413]+z[1413]);
assign {c[1415],s[1414]} = (x[1414]+y[1414]+z[1414]);
assign {c[1416],s[1415]} = (x[1415]+y[1415]+z[1415]);
assign {c[1417],s[1416]} = (x[1416]+y[1416]+z[1416]);
assign {c[1418],s[1417]} = (x[1417]+y[1417]+z[1417]);
assign {c[1419],s[1418]} = (x[1418]+y[1418]+z[1418]);
assign {c[1420],s[1419]} = (x[1419]+y[1419]+z[1419]);
assign {c[1421],s[1420]} = (x[1420]+y[1420]+z[1420]);
assign {c[1422],s[1421]} = (x[1421]+y[1421]+z[1421]);
assign {c[1423],s[1422]} = (x[1422]+y[1422]+z[1422]);
assign {c[1424],s[1423]} = (x[1423]+y[1423]+z[1423]);
assign {c[1425],s[1424]} = (x[1424]+y[1424]+z[1424]);
assign {c[1426],s[1425]} = (x[1425]+y[1425]+z[1425]);
assign {c[1427],s[1426]} = (x[1426]+y[1426]+z[1426]);
assign {c[1428],s[1427]} = (x[1427]+y[1427]+z[1427]);
assign {c[1429],s[1428]} = (x[1428]+y[1428]+z[1428]);
assign {c[1430],s[1429]} = (x[1429]+y[1429]+z[1429]);
assign {c[1431],s[1430]} = (x[1430]+y[1430]+z[1430]);
assign {c[1432],s[1431]} = (x[1431]+y[1431]+z[1431]);
assign {c[1433],s[1432]} = (x[1432]+y[1432]+z[1432]);
assign {c[1434],s[1433]} = (x[1433]+y[1433]+z[1433]);
assign {c[1435],s[1434]} = (x[1434]+y[1434]+z[1434]);
assign {c[1436],s[1435]} = (x[1435]+y[1435]+z[1435]);
assign {c[1437],s[1436]} = (x[1436]+y[1436]+z[1436]);
assign {c[1438],s[1437]} = (x[1437]+y[1437]+z[1437]);
assign {c[1439],s[1438]} = (x[1438]+y[1438]+z[1438]);
assign {c[1440],s[1439]} = (x[1439]+y[1439]+z[1439]);
assign {c[1441],s[1440]} = (x[1440]+y[1440]+z[1440]);
assign {c[1442],s[1441]} = (x[1441]+y[1441]+z[1441]);
assign {c[1443],s[1442]} = (x[1442]+y[1442]+z[1442]);
assign {c[1444],s[1443]} = (x[1443]+y[1443]+z[1443]);
assign {c[1445],s[1444]} = (x[1444]+y[1444]+z[1444]);
assign {c[1446],s[1445]} = (x[1445]+y[1445]+z[1445]);
assign {c[1447],s[1446]} = (x[1446]+y[1446]+z[1446]);
assign {c[1448],s[1447]} = (x[1447]+y[1447]+z[1447]);
assign {c[1449],s[1448]} = (x[1448]+y[1448]+z[1448]);
assign {c[1450],s[1449]} = (x[1449]+y[1449]+z[1449]);
assign {c[1451],s[1450]} = (x[1450]+y[1450]+z[1450]);
assign {c[1452],s[1451]} = (x[1451]+y[1451]+z[1451]);
assign {c[1453],s[1452]} = (x[1452]+y[1452]+z[1452]);
assign {c[1454],s[1453]} = (x[1453]+y[1453]+z[1453]);
assign {c[1455],s[1454]} = (x[1454]+y[1454]+z[1454]);
assign {c[1456],s[1455]} = (x[1455]+y[1455]+z[1455]);
assign {c[1457],s[1456]} = (x[1456]+y[1456]+z[1456]);
assign {c[1458],s[1457]} = (x[1457]+y[1457]+z[1457]);
assign {c[1459],s[1458]} = (x[1458]+y[1458]+z[1458]);
assign {c[1460],s[1459]} = (x[1459]+y[1459]+z[1459]);
assign {c[1461],s[1460]} = (x[1460]+y[1460]+z[1460]);
assign {c[1462],s[1461]} = (x[1461]+y[1461]+z[1461]);
assign {c[1463],s[1462]} = (x[1462]+y[1462]+z[1462]);
assign {c[1464],s[1463]} = (x[1463]+y[1463]+z[1463]);
assign {c[1465],s[1464]} = (x[1464]+y[1464]+z[1464]);
assign {c[1466],s[1465]} = (x[1465]+y[1465]+z[1465]);
assign {c[1467],s[1466]} = (x[1466]+y[1466]+z[1466]);
assign {c[1468],s[1467]} = (x[1467]+y[1467]+z[1467]);
assign {c[1469],s[1468]} = (x[1468]+y[1468]+z[1468]);
assign {c[1470],s[1469]} = (x[1469]+y[1469]+z[1469]);
assign {c[1471],s[1470]} = (x[1470]+y[1470]+z[1470]);
assign {c[1472],s[1471]} = (x[1471]+y[1471]+z[1471]);
assign {c[1473],s[1472]} = (x[1472]+y[1472]+z[1472]);
assign {c[1474],s[1473]} = (x[1473]+y[1473]+z[1473]);
assign {c[1475],s[1474]} = (x[1474]+y[1474]+z[1474]);
assign {c[1476],s[1475]} = (x[1475]+y[1475]+z[1475]);
assign {c[1477],s[1476]} = (x[1476]+y[1476]+z[1476]);
assign {c[1478],s[1477]} = (x[1477]+y[1477]+z[1477]);
assign {c[1479],s[1478]} = (x[1478]+y[1478]+z[1478]);
assign {c[1480],s[1479]} = (x[1479]+y[1479]+z[1479]);
assign {c[1481],s[1480]} = (x[1480]+y[1480]+z[1480]);
assign {c[1482],s[1481]} = (x[1481]+y[1481]+z[1481]);
assign {c[1483],s[1482]} = (x[1482]+y[1482]+z[1482]);
assign {c[1484],s[1483]} = (x[1483]+y[1483]+z[1483]);
assign {c[1485],s[1484]} = (x[1484]+y[1484]+z[1484]);
assign {c[1486],s[1485]} = (x[1485]+y[1485]+z[1485]);
assign {c[1487],s[1486]} = (x[1486]+y[1486]+z[1486]);
assign {c[1488],s[1487]} = (x[1487]+y[1487]+z[1487]);
assign {c[1489],s[1488]} = (x[1488]+y[1488]+z[1488]);
assign {c[1490],s[1489]} = (x[1489]+y[1489]+z[1489]);
assign {c[1491],s[1490]} = (x[1490]+y[1490]+z[1490]);
assign {c[1492],s[1491]} = (x[1491]+y[1491]+z[1491]);
assign {c[1493],s[1492]} = (x[1492]+y[1492]+z[1492]);
assign {c[1494],s[1493]} = (x[1493]+y[1493]+z[1493]);
assign {c[1495],s[1494]} = (x[1494]+y[1494]+z[1494]);
assign {c[1496],s[1495]} = (x[1495]+y[1495]+z[1495]);
assign {c[1497],s[1496]} = (x[1496]+y[1496]+z[1496]);
assign {c[1498],s[1497]} = (x[1497]+y[1497]+z[1497]);
assign {c[1499],s[1498]} = (x[1498]+y[1498]+z[1498]);
assign {c[1500],s[1499]} = (x[1499]+y[1499]+z[1499]);
assign {c[1501],s[1500]} = (x[1500]+y[1500]+z[1500]);
assign {c[1502],s[1501]} = (x[1501]+y[1501]+z[1501]);
assign {c[1503],s[1502]} = (x[1502]+y[1502]+z[1502]);
assign {c[1504],s[1503]} = (x[1503]+y[1503]+z[1503]);
assign {c[1505],s[1504]} = (x[1504]+y[1504]+z[1504]);
assign {c[1506],s[1505]} = (x[1505]+y[1505]+z[1505]);
assign {c[1507],s[1506]} = (x[1506]+y[1506]+z[1506]);
assign {c[1508],s[1507]} = (x[1507]+y[1507]+z[1507]);
assign {c[1509],s[1508]} = (x[1508]+y[1508]+z[1508]);
assign {c[1510],s[1509]} = (x[1509]+y[1509]+z[1509]);
assign {c[1511],s[1510]} = (x[1510]+y[1510]+z[1510]);
assign {c[1512],s[1511]} = (x[1511]+y[1511]+z[1511]);
assign {c[1513],s[1512]} = (x[1512]+y[1512]+z[1512]);
assign {c[1514],s[1513]} = (x[1513]+y[1513]+z[1513]);
assign {c[1515],s[1514]} = (x[1514]+y[1514]+z[1514]);
assign {c[1516],s[1515]} = (x[1515]+y[1515]+z[1515]);
assign {c[1517],s[1516]} = (x[1516]+y[1516]+z[1516]);
assign {c[1518],s[1517]} = (x[1517]+y[1517]+z[1517]);
assign {c[1519],s[1518]} = (x[1518]+y[1518]+z[1518]);
assign {c[1520],s[1519]} = (x[1519]+y[1519]+z[1519]);
assign {c[1521],s[1520]} = (x[1520]+y[1520]+z[1520]);
assign {c[1522],s[1521]} = (x[1521]+y[1521]+z[1521]);
assign {c[1523],s[1522]} = (x[1522]+y[1522]+z[1522]);
assign {c[1524],s[1523]} = (x[1523]+y[1523]+z[1523]);
assign {c[1525],s[1524]} = (x[1524]+y[1524]+z[1524]);
assign {c[1526],s[1525]} = (x[1525]+y[1525]+z[1525]);
assign {c[1527],s[1526]} = (x[1526]+y[1526]+z[1526]);
assign {c[1528],s[1527]} = (x[1527]+y[1527]+z[1527]);
assign {c[1529],s[1528]} = (x[1528]+y[1528]+z[1528]);
assign {c[1530],s[1529]} = (x[1529]+y[1529]+z[1529]);
assign {c[1531],s[1530]} = (x[1530]+y[1530]+z[1530]);
assign {c[1532],s[1531]} = (x[1531]+y[1531]+z[1531]);
assign {c[1533],s[1532]} = (x[1532]+y[1532]+z[1532]);
assign {c[1534],s[1533]} = (x[1533]+y[1533]+z[1533]);
assign {c[1535],s[1534]} = (x[1534]+y[1534]+z[1534]);
assign {c[1536],s[1535]} = (x[1535]+y[1535]+z[1535]);
assign {c[1537],s[1536]} = (x[1536]+y[1536]+z[1536]);
assign {c[1538],s[1537]} = (x[1537]+y[1537]+z[1537]);
assign {c[1539],s[1538]} = (x[1538]+y[1538]+z[1538]);
assign {c[1540],s[1539]} = (x[1539]+y[1539]+z[1539]);
assign {c[1541],s[1540]} = (x[1540]+y[1540]+z[1540]);
assign {c[1542],s[1541]} = (x[1541]+y[1541]+z[1541]);
assign {c[1543],s[1542]} = (x[1542]+y[1542]+z[1542]);
assign {c[1544],s[1543]} = (x[1543]+y[1543]+z[1543]);
assign {c[1545],s[1544]} = (x[1544]+y[1544]+z[1544]);
assign {c[1546],s[1545]} = (x[1545]+y[1545]+z[1545]);
assign {c[1547],s[1546]} = (x[1546]+y[1546]+z[1546]);
assign {c[1548],s[1547]} = (x[1547]+y[1547]+z[1547]);
assign {c[1549],s[1548]} = (x[1548]+y[1548]+z[1548]);
assign {c[1550],s[1549]} = (x[1549]+y[1549]+z[1549]);
assign {c[1551],s[1550]} = (x[1550]+y[1550]+z[1550]);
assign {c[1552],s[1551]} = (x[1551]+y[1551]+z[1551]);
assign {c[1553],s[1552]} = (x[1552]+y[1552]+z[1552]);
assign {c[1554],s[1553]} = (x[1553]+y[1553]+z[1553]);
assign {c[1555],s[1554]} = (x[1554]+y[1554]+z[1554]);
assign {c[1556],s[1555]} = (x[1555]+y[1555]+z[1555]);
assign {c[1557],s[1556]} = (x[1556]+y[1556]+z[1556]);
assign {c[1558],s[1557]} = (x[1557]+y[1557]+z[1557]);
assign {c[1559],s[1558]} = (x[1558]+y[1558]+z[1558]);
assign {c[1560],s[1559]} = (x[1559]+y[1559]+z[1559]);
assign {c[1561],s[1560]} = (x[1560]+y[1560]+z[1560]);
assign {c[1562],s[1561]} = (x[1561]+y[1561]+z[1561]);
assign {c[1563],s[1562]} = (x[1562]+y[1562]+z[1562]);
assign {c[1564],s[1563]} = (x[1563]+y[1563]+z[1563]);
assign {c[1565],s[1564]} = (x[1564]+y[1564]+z[1564]);
assign {c[1566],s[1565]} = (x[1565]+y[1565]+z[1565]);
assign {c[1567],s[1566]} = (x[1566]+y[1566]+z[1566]);
assign {c[1568],s[1567]} = (x[1567]+y[1567]+z[1567]);
assign {c[1569],s[1568]} = (x[1568]+y[1568]+z[1568]);
assign {c[1570],s[1569]} = (x[1569]+y[1569]+z[1569]);
assign {c[1571],s[1570]} = (x[1570]+y[1570]+z[1570]);
assign {c[1572],s[1571]} = (x[1571]+y[1571]+z[1571]);
assign {c[1573],s[1572]} = (x[1572]+y[1572]+z[1572]);
assign {c[1574],s[1573]} = (x[1573]+y[1573]+z[1573]);
assign {c[1575],s[1574]} = (x[1574]+y[1574]+z[1574]);
assign {c[1576],s[1575]} = (x[1575]+y[1575]+z[1575]);
assign {c[1577],s[1576]} = (x[1576]+y[1576]+z[1576]);
assign {c[1578],s[1577]} = (x[1577]+y[1577]+z[1577]);
assign {c[1579],s[1578]} = (x[1578]+y[1578]+z[1578]);
assign {c[1580],s[1579]} = (x[1579]+y[1579]+z[1579]);
assign {c[1581],s[1580]} = (x[1580]+y[1580]+z[1580]);
assign {c[1582],s[1581]} = (x[1581]+y[1581]+z[1581]);
assign {c[1583],s[1582]} = (x[1582]+y[1582]+z[1582]);
assign {c[1584],s[1583]} = (x[1583]+y[1583]+z[1583]);
assign {c[1585],s[1584]} = (x[1584]+y[1584]+z[1584]);
assign {c[1586],s[1585]} = (x[1585]+y[1585]+z[1585]);
assign {c[1587],s[1586]} = (x[1586]+y[1586]+z[1586]);
assign {c[1588],s[1587]} = (x[1587]+y[1587]+z[1587]);
assign {c[1589],s[1588]} = (x[1588]+y[1588]+z[1588]);
assign {c[1590],s[1589]} = (x[1589]+y[1589]+z[1589]);
assign {c[1591],s[1590]} = (x[1590]+y[1590]+z[1590]);
assign {c[1592],s[1591]} = (x[1591]+y[1591]+z[1591]);
assign {c[1593],s[1592]} = (x[1592]+y[1592]+z[1592]);
assign {c[1594],s[1593]} = (x[1593]+y[1593]+z[1593]);
assign {c[1595],s[1594]} = (x[1594]+y[1594]+z[1594]);
assign {c[1596],s[1595]} = (x[1595]+y[1595]+z[1595]);
assign {c[1597],s[1596]} = (x[1596]+y[1596]+z[1596]);
assign {c[1598],s[1597]} = (x[1597]+y[1597]+z[1597]);
assign {c[1599],s[1598]} = (x[1598]+y[1598]+z[1598]);
assign {c[1600],s[1599]} = (x[1599]+y[1599]+z[1599]);
assign {c[1601],s[1600]} = (x[1600]+y[1600]+z[1600]);
assign {c[1602],s[1601]} = (x[1601]+y[1601]+z[1601]);
assign {c[1603],s[1602]} = (x[1602]+y[1602]+z[1602]);
assign {c[1604],s[1603]} = (x[1603]+y[1603]+z[1603]);
assign {c[1605],s[1604]} = (x[1604]+y[1604]+z[1604]);
assign {c[1606],s[1605]} = (x[1605]+y[1605]+z[1605]);
assign {c[1607],s[1606]} = (x[1606]+y[1606]+z[1606]);
assign {c[1608],s[1607]} = (x[1607]+y[1607]+z[1607]);
assign {c[1609],s[1608]} = (x[1608]+y[1608]+z[1608]);
assign {c[1610],s[1609]} = (x[1609]+y[1609]+z[1609]);
assign {c[1611],s[1610]} = (x[1610]+y[1610]+z[1610]);
assign {c[1612],s[1611]} = (x[1611]+y[1611]+z[1611]);
assign {c[1613],s[1612]} = (x[1612]+y[1612]+z[1612]);
assign {c[1614],s[1613]} = (x[1613]+y[1613]+z[1613]);
assign {c[1615],s[1614]} = (x[1614]+y[1614]+z[1614]);
assign {c[1616],s[1615]} = (x[1615]+y[1615]+z[1615]);
assign {c[1617],s[1616]} = (x[1616]+y[1616]+z[1616]);
assign {c[1618],s[1617]} = (x[1617]+y[1617]+z[1617]);
assign {c[1619],s[1618]} = (x[1618]+y[1618]+z[1618]);
assign {c[1620],s[1619]} = (x[1619]+y[1619]+z[1619]);
assign {c[1621],s[1620]} = (x[1620]+y[1620]+z[1620]);
assign {c[1622],s[1621]} = (x[1621]+y[1621]+z[1621]);
assign {c[1623],s[1622]} = (x[1622]+y[1622]+z[1622]);
assign {c[1624],s[1623]} = (x[1623]+y[1623]+z[1623]);
assign {c[1625],s[1624]} = (x[1624]+y[1624]+z[1624]);
assign {c[1626],s[1625]} = (x[1625]+y[1625]+z[1625]);
assign {c[1627],s[1626]} = (x[1626]+y[1626]+z[1626]);
assign {c[1628],s[1627]} = (x[1627]+y[1627]+z[1627]);
assign {c[1629],s[1628]} = (x[1628]+y[1628]+z[1628]);
assign {c[1630],s[1629]} = (x[1629]+y[1629]+z[1629]);
assign {c[1631],s[1630]} = (x[1630]+y[1630]+z[1630]);
assign {c[1632],s[1631]} = (x[1631]+y[1631]+z[1631]);
assign {c[1633],s[1632]} = (x[1632]+y[1632]+z[1632]);
assign {c[1634],s[1633]} = (x[1633]+y[1633]+z[1633]);
assign {c[1635],s[1634]} = (x[1634]+y[1634]+z[1634]);
assign {c[1636],s[1635]} = (x[1635]+y[1635]+z[1635]);
assign {c[1637],s[1636]} = (x[1636]+y[1636]+z[1636]);
assign {c[1638],s[1637]} = (x[1637]+y[1637]+z[1637]);
assign {c[1639],s[1638]} = (x[1638]+y[1638]+z[1638]);
assign {c[1640],s[1639]} = (x[1639]+y[1639]+z[1639]);
assign {c[1641],s[1640]} = (x[1640]+y[1640]+z[1640]);
assign {c[1642],s[1641]} = (x[1641]+y[1641]+z[1641]);
assign {c[1643],s[1642]} = (x[1642]+y[1642]+z[1642]);
assign {c[1644],s[1643]} = (x[1643]+y[1643]+z[1643]);
assign {c[1645],s[1644]} = (x[1644]+y[1644]+z[1644]);
assign {c[1646],s[1645]} = (x[1645]+y[1645]+z[1645]);
assign {c[1647],s[1646]} = (x[1646]+y[1646]+z[1646]);
assign {c[1648],s[1647]} = (x[1647]+y[1647]+z[1647]);
assign {c[1649],s[1648]} = (x[1648]+y[1648]+z[1648]);
assign {c[1650],s[1649]} = (x[1649]+y[1649]+z[1649]);
assign {c[1651],s[1650]} = (x[1650]+y[1650]+z[1650]);
assign {c[1652],s[1651]} = (x[1651]+y[1651]+z[1651]);
assign {c[1653],s[1652]} = (x[1652]+y[1652]+z[1652]);
assign {c[1654],s[1653]} = (x[1653]+y[1653]+z[1653]);
assign {c[1655],s[1654]} = (x[1654]+y[1654]+z[1654]);
assign {c[1656],s[1655]} = (x[1655]+y[1655]+z[1655]);
assign {c[1657],s[1656]} = (x[1656]+y[1656]+z[1656]);
assign {c[1658],s[1657]} = (x[1657]+y[1657]+z[1657]);
assign {c[1659],s[1658]} = (x[1658]+y[1658]+z[1658]);
assign {c[1660],s[1659]} = (x[1659]+y[1659]+z[1659]);
assign {c[1661],s[1660]} = (x[1660]+y[1660]+z[1660]);
assign {c[1662],s[1661]} = (x[1661]+y[1661]+z[1661]);
assign {c[1663],s[1662]} = (x[1662]+y[1662]+z[1662]);
assign {c[1664],s[1663]} = (x[1663]+y[1663]+z[1663]);
assign {c[1665],s[1664]} = (x[1664]+y[1664]+z[1664]);
assign {c[1666],s[1665]} = (x[1665]+y[1665]+z[1665]);
assign {c[1667],s[1666]} = (x[1666]+y[1666]+z[1666]);
assign {c[1668],s[1667]} = (x[1667]+y[1667]+z[1667]);
assign {c[1669],s[1668]} = (x[1668]+y[1668]+z[1668]);
assign {c[1670],s[1669]} = (x[1669]+y[1669]+z[1669]);
assign {c[1671],s[1670]} = (x[1670]+y[1670]+z[1670]);
assign {c[1672],s[1671]} = (x[1671]+y[1671]+z[1671]);
assign {c[1673],s[1672]} = (x[1672]+y[1672]+z[1672]);
assign {c[1674],s[1673]} = (x[1673]+y[1673]+z[1673]);
assign {c[1675],s[1674]} = (x[1674]+y[1674]+z[1674]);
assign {c[1676],s[1675]} = (x[1675]+y[1675]+z[1675]);
assign {c[1677],s[1676]} = (x[1676]+y[1676]+z[1676]);
assign {c[1678],s[1677]} = (x[1677]+y[1677]+z[1677]);
assign {c[1679],s[1678]} = (x[1678]+y[1678]+z[1678]);
assign {c[1680],s[1679]} = (x[1679]+y[1679]+z[1679]);
assign {c[1681],s[1680]} = (x[1680]+y[1680]+z[1680]);
assign {c[1682],s[1681]} = (x[1681]+y[1681]+z[1681]);
assign {c[1683],s[1682]} = (x[1682]+y[1682]+z[1682]);
assign {c[1684],s[1683]} = (x[1683]+y[1683]+z[1683]);
assign {c[1685],s[1684]} = (x[1684]+y[1684]+z[1684]);
assign {c[1686],s[1685]} = (x[1685]+y[1685]+z[1685]);
assign {c[1687],s[1686]} = (x[1686]+y[1686]+z[1686]);
assign {c[1688],s[1687]} = (x[1687]+y[1687]+z[1687]);
assign {c[1689],s[1688]} = (x[1688]+y[1688]+z[1688]);
assign {c[1690],s[1689]} = (x[1689]+y[1689]+z[1689]);
assign {c[1691],s[1690]} = (x[1690]+y[1690]+z[1690]);
assign {c[1692],s[1691]} = (x[1691]+y[1691]+z[1691]);
assign {c[1693],s[1692]} = (x[1692]+y[1692]+z[1692]);
assign {c[1694],s[1693]} = (x[1693]+y[1693]+z[1693]);
assign {c[1695],s[1694]} = (x[1694]+y[1694]+z[1694]);
assign {c[1696],s[1695]} = (x[1695]+y[1695]+z[1695]);
assign {c[1697],s[1696]} = (x[1696]+y[1696]+z[1696]);
assign {c[1698],s[1697]} = (x[1697]+y[1697]+z[1697]);
assign {c[1699],s[1698]} = (x[1698]+y[1698]+z[1698]);
assign {c[1700],s[1699]} = (x[1699]+y[1699]+z[1699]);
assign {c[1701],s[1700]} = (x[1700]+y[1700]+z[1700]);
assign {c[1702],s[1701]} = (x[1701]+y[1701]+z[1701]);
assign {c[1703],s[1702]} = (x[1702]+y[1702]+z[1702]);
assign {c[1704],s[1703]} = (x[1703]+y[1703]+z[1703]);
assign {c[1705],s[1704]} = (x[1704]+y[1704]+z[1704]);
assign {c[1706],s[1705]} = (x[1705]+y[1705]+z[1705]);
assign {c[1707],s[1706]} = (x[1706]+y[1706]+z[1706]);
assign {c[1708],s[1707]} = (x[1707]+y[1707]+z[1707]);
assign {c[1709],s[1708]} = (x[1708]+y[1708]+z[1708]);
assign {c[1710],s[1709]} = (x[1709]+y[1709]+z[1709]);
assign {c[1711],s[1710]} = (x[1710]+y[1710]+z[1710]);
assign {c[1712],s[1711]} = (x[1711]+y[1711]+z[1711]);
assign {c[1713],s[1712]} = (x[1712]+y[1712]+z[1712]);
assign {c[1714],s[1713]} = (x[1713]+y[1713]+z[1713]);
assign {c[1715],s[1714]} = (x[1714]+y[1714]+z[1714]);
assign {c[1716],s[1715]} = (x[1715]+y[1715]+z[1715]);
assign {c[1717],s[1716]} = (x[1716]+y[1716]+z[1716]);
assign {c[1718],s[1717]} = (x[1717]+y[1717]+z[1717]);
assign {c[1719],s[1718]} = (x[1718]+y[1718]+z[1718]);
assign {c[1720],s[1719]} = (x[1719]+y[1719]+z[1719]);
assign {c[1721],s[1720]} = (x[1720]+y[1720]+z[1720]);
assign {c[1722],s[1721]} = (x[1721]+y[1721]+z[1721]);
assign {c[1723],s[1722]} = (x[1722]+y[1722]+z[1722]);
assign {c[1724],s[1723]} = (x[1723]+y[1723]+z[1723]);
assign {c[1725],s[1724]} = (x[1724]+y[1724]+z[1724]);
assign {c[1726],s[1725]} = (x[1725]+y[1725]+z[1725]);
assign {c[1727],s[1726]} = (x[1726]+y[1726]+z[1726]);
assign {c[1728],s[1727]} = (x[1727]+y[1727]+z[1727]);
assign {c[1729],s[1728]} = (x[1728]+y[1728]+z[1728]);
assign {c[1730],s[1729]} = (x[1729]+y[1729]+z[1729]);
assign {c[1731],s[1730]} = (x[1730]+y[1730]+z[1730]);
assign {c[1732],s[1731]} = (x[1731]+y[1731]+z[1731]);
assign {c[1733],s[1732]} = (x[1732]+y[1732]+z[1732]);
assign {c[1734],s[1733]} = (x[1733]+y[1733]+z[1733]);
assign {c[1735],s[1734]} = (x[1734]+y[1734]+z[1734]);
assign {c[1736],s[1735]} = (x[1735]+y[1735]+z[1735]);
assign {c[1737],s[1736]} = (x[1736]+y[1736]+z[1736]);
assign {c[1738],s[1737]} = (x[1737]+y[1737]+z[1737]);
assign {c[1739],s[1738]} = (x[1738]+y[1738]+z[1738]);
assign {c[1740],s[1739]} = (x[1739]+y[1739]+z[1739]);
assign {c[1741],s[1740]} = (x[1740]+y[1740]+z[1740]);
assign {c[1742],s[1741]} = (x[1741]+y[1741]+z[1741]);
assign {c[1743],s[1742]} = (x[1742]+y[1742]+z[1742]);
assign {c[1744],s[1743]} = (x[1743]+y[1743]+z[1743]);
assign {c[1745],s[1744]} = (x[1744]+y[1744]+z[1744]);
assign {c[1746],s[1745]} = (x[1745]+y[1745]+z[1745]);
assign {c[1747],s[1746]} = (x[1746]+y[1746]+z[1746]);
assign {c[1748],s[1747]} = (x[1747]+y[1747]+z[1747]);
assign {c[1749],s[1748]} = (x[1748]+y[1748]+z[1748]);
assign {c[1750],s[1749]} = (x[1749]+y[1749]+z[1749]);
assign {c[1751],s[1750]} = (x[1750]+y[1750]+z[1750]);
assign {c[1752],s[1751]} = (x[1751]+y[1751]+z[1751]);
assign {c[1753],s[1752]} = (x[1752]+y[1752]+z[1752]);
assign {c[1754],s[1753]} = (x[1753]+y[1753]+z[1753]);
assign {c[1755],s[1754]} = (x[1754]+y[1754]+z[1754]);
assign {c[1756],s[1755]} = (x[1755]+y[1755]+z[1755]);
assign {c[1757],s[1756]} = (x[1756]+y[1756]+z[1756]);
assign {c[1758],s[1757]} = (x[1757]+y[1757]+z[1757]);
assign {c[1759],s[1758]} = (x[1758]+y[1758]+z[1758]);
assign {c[1760],s[1759]} = (x[1759]+y[1759]+z[1759]);
assign {c[1761],s[1760]} = (x[1760]+y[1760]+z[1760]);
assign {c[1762],s[1761]} = (x[1761]+y[1761]+z[1761]);
assign {c[1763],s[1762]} = (x[1762]+y[1762]+z[1762]);
assign {c[1764],s[1763]} = (x[1763]+y[1763]+z[1763]);
assign {c[1765],s[1764]} = (x[1764]+y[1764]+z[1764]);
assign {c[1766],s[1765]} = (x[1765]+y[1765]+z[1765]);
assign {c[1767],s[1766]} = (x[1766]+y[1766]+z[1766]);
assign {c[1768],s[1767]} = (x[1767]+y[1767]+z[1767]);
assign {c[1769],s[1768]} = (x[1768]+y[1768]+z[1768]);
assign {c[1770],s[1769]} = (x[1769]+y[1769]+z[1769]);
assign {c[1771],s[1770]} = (x[1770]+y[1770]+z[1770]);
assign {c[1772],s[1771]} = (x[1771]+y[1771]+z[1771]);
assign {c[1773],s[1772]} = (x[1772]+y[1772]+z[1772]);
assign {c[1774],s[1773]} = (x[1773]+y[1773]+z[1773]);
assign {c[1775],s[1774]} = (x[1774]+y[1774]+z[1774]);
assign {c[1776],s[1775]} = (x[1775]+y[1775]+z[1775]);
assign {c[1777],s[1776]} = (x[1776]+y[1776]+z[1776]);
assign {c[1778],s[1777]} = (x[1777]+y[1777]+z[1777]);
assign {c[1779],s[1778]} = (x[1778]+y[1778]+z[1778]);
assign {c[1780],s[1779]} = (x[1779]+y[1779]+z[1779]);
assign {c[1781],s[1780]} = (x[1780]+y[1780]+z[1780]);
assign {c[1782],s[1781]} = (x[1781]+y[1781]+z[1781]);
assign {c[1783],s[1782]} = (x[1782]+y[1782]+z[1782]);
assign {c[1784],s[1783]} = (x[1783]+y[1783]+z[1783]);
assign {c[1785],s[1784]} = (x[1784]+y[1784]+z[1784]);
assign {c[1786],s[1785]} = (x[1785]+y[1785]+z[1785]);
assign {c[1787],s[1786]} = (x[1786]+y[1786]+z[1786]);
assign {c[1788],s[1787]} = (x[1787]+y[1787]+z[1787]);
assign {c[1789],s[1788]} = (x[1788]+y[1788]+z[1788]);
assign {c[1790],s[1789]} = (x[1789]+y[1789]+z[1789]);
assign {c[1791],s[1790]} = (x[1790]+y[1790]+z[1790]);
assign {c[1792],s[1791]} = (x[1791]+y[1791]+z[1791]);
assign {c[1793],s[1792]} = (x[1792]+y[1792]+z[1792]);
assign {c[1794],s[1793]} = (x[1793]+y[1793]+z[1793]);
assign {c[1795],s[1794]} = (x[1794]+y[1794]+z[1794]);
assign {c[1796],s[1795]} = (x[1795]+y[1795]+z[1795]);
assign {c[1797],s[1796]} = (x[1796]+y[1796]+z[1796]);
assign {c[1798],s[1797]} = (x[1797]+y[1797]+z[1797]);
assign {c[1799],s[1798]} = (x[1798]+y[1798]+z[1798]);
assign {c[1800],s[1799]} = (x[1799]+y[1799]+z[1799]);
assign {c[1801],s[1800]} = (x[1800]+y[1800]+z[1800]);
assign {c[1802],s[1801]} = (x[1801]+y[1801]+z[1801]);
assign {c[1803],s[1802]} = (x[1802]+y[1802]+z[1802]);
assign {c[1804],s[1803]} = (x[1803]+y[1803]+z[1803]);
assign {c[1805],s[1804]} = (x[1804]+y[1804]+z[1804]);
assign {c[1806],s[1805]} = (x[1805]+y[1805]+z[1805]);
assign {c[1807],s[1806]} = (x[1806]+y[1806]+z[1806]);
assign {c[1808],s[1807]} = (x[1807]+y[1807]+z[1807]);
assign {c[1809],s[1808]} = (x[1808]+y[1808]+z[1808]);
assign {c[1810],s[1809]} = (x[1809]+y[1809]+z[1809]);
assign {c[1811],s[1810]} = (x[1810]+y[1810]+z[1810]);
assign {c[1812],s[1811]} = (x[1811]+y[1811]+z[1811]);
assign {c[1813],s[1812]} = (x[1812]+y[1812]+z[1812]);
assign {c[1814],s[1813]} = (x[1813]+y[1813]+z[1813]);
assign {c[1815],s[1814]} = (x[1814]+y[1814]+z[1814]);
assign {c[1816],s[1815]} = (x[1815]+y[1815]+z[1815]);
assign {c[1817],s[1816]} = (x[1816]+y[1816]+z[1816]);
assign {c[1818],s[1817]} = (x[1817]+y[1817]+z[1817]);
assign {c[1819],s[1818]} = (x[1818]+y[1818]+z[1818]);
assign {c[1820],s[1819]} = (x[1819]+y[1819]+z[1819]);
assign {c[1821],s[1820]} = (x[1820]+y[1820]+z[1820]);
assign {c[1822],s[1821]} = (x[1821]+y[1821]+z[1821]);
assign {c[1823],s[1822]} = (x[1822]+y[1822]+z[1822]);
assign {c[1824],s[1823]} = (x[1823]+y[1823]+z[1823]);
assign {c[1825],s[1824]} = (x[1824]+y[1824]+z[1824]);
assign {c[1826],s[1825]} = (x[1825]+y[1825]+z[1825]);
assign {c[1827],s[1826]} = (x[1826]+y[1826]+z[1826]);
assign {c[1828],s[1827]} = (x[1827]+y[1827]+z[1827]);
assign {c[1829],s[1828]} = (x[1828]+y[1828]+z[1828]);
assign {c[1830],s[1829]} = (x[1829]+y[1829]+z[1829]);
assign {c[1831],s[1830]} = (x[1830]+y[1830]+z[1830]);
assign {c[1832],s[1831]} = (x[1831]+y[1831]+z[1831]);
assign {c[1833],s[1832]} = (x[1832]+y[1832]+z[1832]);
assign {c[1834],s[1833]} = (x[1833]+y[1833]+z[1833]);
assign {c[1835],s[1834]} = (x[1834]+y[1834]+z[1834]);
assign {c[1836],s[1835]} = (x[1835]+y[1835]+z[1835]);
assign {c[1837],s[1836]} = (x[1836]+y[1836]+z[1836]);
assign {c[1838],s[1837]} = (x[1837]+y[1837]+z[1837]);
assign {c[1839],s[1838]} = (x[1838]+y[1838]+z[1838]);
assign {c[1840],s[1839]} = (x[1839]+y[1839]+z[1839]);
assign {c[1841],s[1840]} = (x[1840]+y[1840]+z[1840]);
assign {c[1842],s[1841]} = (x[1841]+y[1841]+z[1841]);
assign {c[1843],s[1842]} = (x[1842]+y[1842]+z[1842]);
assign {c[1844],s[1843]} = (x[1843]+y[1843]+z[1843]);
assign {c[1845],s[1844]} = (x[1844]+y[1844]+z[1844]);
assign {c[1846],s[1845]} = (x[1845]+y[1845]+z[1845]);
assign {c[1847],s[1846]} = (x[1846]+y[1846]+z[1846]);
assign {c[1848],s[1847]} = (x[1847]+y[1847]+z[1847]);
assign {c[1849],s[1848]} = (x[1848]+y[1848]+z[1848]);
assign {c[1850],s[1849]} = (x[1849]+y[1849]+z[1849]);
assign {c[1851],s[1850]} = (x[1850]+y[1850]+z[1850]);
assign {c[1852],s[1851]} = (x[1851]+y[1851]+z[1851]);
assign {c[1853],s[1852]} = (x[1852]+y[1852]+z[1852]);
assign {c[1854],s[1853]} = (x[1853]+y[1853]+z[1853]);
assign {c[1855],s[1854]} = (x[1854]+y[1854]+z[1854]);
assign {c[1856],s[1855]} = (x[1855]+y[1855]+z[1855]);
assign {c[1857],s[1856]} = (x[1856]+y[1856]+z[1856]);
assign {c[1858],s[1857]} = (x[1857]+y[1857]+z[1857]);
assign {c[1859],s[1858]} = (x[1858]+y[1858]+z[1858]);
assign {c[1860],s[1859]} = (x[1859]+y[1859]+z[1859]);
assign {c[1861],s[1860]} = (x[1860]+y[1860]+z[1860]);
assign {c[1862],s[1861]} = (x[1861]+y[1861]+z[1861]);
assign {c[1863],s[1862]} = (x[1862]+y[1862]+z[1862]);
assign {c[1864],s[1863]} = (x[1863]+y[1863]+z[1863]);
assign {c[1865],s[1864]} = (x[1864]+y[1864]+z[1864]);
assign {c[1866],s[1865]} = (x[1865]+y[1865]+z[1865]);
assign {c[1867],s[1866]} = (x[1866]+y[1866]+z[1866]);
assign {c[1868],s[1867]} = (x[1867]+y[1867]+z[1867]);
assign {c[1869],s[1868]} = (x[1868]+y[1868]+z[1868]);
assign {c[1870],s[1869]} = (x[1869]+y[1869]+z[1869]);
assign {c[1871],s[1870]} = (x[1870]+y[1870]+z[1870]);
assign {c[1872],s[1871]} = (x[1871]+y[1871]+z[1871]);
assign {c[1873],s[1872]} = (x[1872]+y[1872]+z[1872]);
assign {c[1874],s[1873]} = (x[1873]+y[1873]+z[1873]);
assign {c[1875],s[1874]} = (x[1874]+y[1874]+z[1874]);
assign {c[1876],s[1875]} = (x[1875]+y[1875]+z[1875]);
assign {c[1877],s[1876]} = (x[1876]+y[1876]+z[1876]);
assign {c[1878],s[1877]} = (x[1877]+y[1877]+z[1877]);
assign {c[1879],s[1878]} = (x[1878]+y[1878]+z[1878]);
assign {c[1880],s[1879]} = (x[1879]+y[1879]+z[1879]);
assign {c[1881],s[1880]} = (x[1880]+y[1880]+z[1880]);
assign {c[1882],s[1881]} = (x[1881]+y[1881]+z[1881]);
assign {c[1883],s[1882]} = (x[1882]+y[1882]+z[1882]);
assign {c[1884],s[1883]} = (x[1883]+y[1883]+z[1883]);
assign {c[1885],s[1884]} = (x[1884]+y[1884]+z[1884]);
assign {c[1886],s[1885]} = (x[1885]+y[1885]+z[1885]);
assign {c[1887],s[1886]} = (x[1886]+y[1886]+z[1886]);
assign {c[1888],s[1887]} = (x[1887]+y[1887]+z[1887]);
assign {c[1889],s[1888]} = (x[1888]+y[1888]+z[1888]);
assign {c[1890],s[1889]} = (x[1889]+y[1889]+z[1889]);
assign {c[1891],s[1890]} = (x[1890]+y[1890]+z[1890]);
assign {c[1892],s[1891]} = (x[1891]+y[1891]+z[1891]);
assign {c[1893],s[1892]} = (x[1892]+y[1892]+z[1892]);
assign {c[1894],s[1893]} = (x[1893]+y[1893]+z[1893]);
assign {c[1895],s[1894]} = (x[1894]+y[1894]+z[1894]);
assign {c[1896],s[1895]} = (x[1895]+y[1895]+z[1895]);
assign {c[1897],s[1896]} = (x[1896]+y[1896]+z[1896]);
assign {c[1898],s[1897]} = (x[1897]+y[1897]+z[1897]);
assign {c[1899],s[1898]} = (x[1898]+y[1898]+z[1898]);
assign {c[1900],s[1899]} = (x[1899]+y[1899]+z[1899]);
assign {c[1901],s[1900]} = (x[1900]+y[1900]+z[1900]);
assign {c[1902],s[1901]} = (x[1901]+y[1901]+z[1901]);
assign {c[1903],s[1902]} = (x[1902]+y[1902]+z[1902]);
assign {c[1904],s[1903]} = (x[1903]+y[1903]+z[1903]);
assign {c[1905],s[1904]} = (x[1904]+y[1904]+z[1904]);
assign {c[1906],s[1905]} = (x[1905]+y[1905]+z[1905]);
assign {c[1907],s[1906]} = (x[1906]+y[1906]+z[1906]);
assign {c[1908],s[1907]} = (x[1907]+y[1907]+z[1907]);
assign {c[1909],s[1908]} = (x[1908]+y[1908]+z[1908]);
assign {c[1910],s[1909]} = (x[1909]+y[1909]+z[1909]);
assign {c[1911],s[1910]} = (x[1910]+y[1910]+z[1910]);
assign {c[1912],s[1911]} = (x[1911]+y[1911]+z[1911]);
assign {c[1913],s[1912]} = (x[1912]+y[1912]+z[1912]);
assign {c[1914],s[1913]} = (x[1913]+y[1913]+z[1913]);
assign {c[1915],s[1914]} = (x[1914]+y[1914]+z[1914]);
assign {c[1916],s[1915]} = (x[1915]+y[1915]+z[1915]);
assign {c[1917],s[1916]} = (x[1916]+y[1916]+z[1916]);
assign {c[1918],s[1917]} = (x[1917]+y[1917]+z[1917]);
assign {c[1919],s[1918]} = (x[1918]+y[1918]+z[1918]);
assign {c[1920],s[1919]} = (x[1919]+y[1919]+z[1919]);
assign {c[1921],s[1920]} = (x[1920]+y[1920]+z[1920]);
assign {c[1922],s[1921]} = (x[1921]+y[1921]+z[1921]);
assign {c[1923],s[1922]} = (x[1922]+y[1922]+z[1922]);
assign {c[1924],s[1923]} = (x[1923]+y[1923]+z[1923]);
assign {c[1925],s[1924]} = (x[1924]+y[1924]+z[1924]);
assign {c[1926],s[1925]} = (x[1925]+y[1925]+z[1925]);
assign {c[1927],s[1926]} = (x[1926]+y[1926]+z[1926]);
assign {c[1928],s[1927]} = (x[1927]+y[1927]+z[1927]);
assign {c[1929],s[1928]} = (x[1928]+y[1928]+z[1928]);
assign {c[1930],s[1929]} = (x[1929]+y[1929]+z[1929]);
assign {c[1931],s[1930]} = (x[1930]+y[1930]+z[1930]);
assign {c[1932],s[1931]} = (x[1931]+y[1931]+z[1931]);
assign {c[1933],s[1932]} = (x[1932]+y[1932]+z[1932]);
assign {c[1934],s[1933]} = (x[1933]+y[1933]+z[1933]);
assign {c[1935],s[1934]} = (x[1934]+y[1934]+z[1934]);
assign {c[1936],s[1935]} = (x[1935]+y[1935]+z[1935]);
assign {c[1937],s[1936]} = (x[1936]+y[1936]+z[1936]);
assign {c[1938],s[1937]} = (x[1937]+y[1937]+z[1937]);
assign {c[1939],s[1938]} = (x[1938]+y[1938]+z[1938]);
assign {c[1940],s[1939]} = (x[1939]+y[1939]+z[1939]);
assign {c[1941],s[1940]} = (x[1940]+y[1940]+z[1940]);
assign {c[1942],s[1941]} = (x[1941]+y[1941]+z[1941]);
assign {c[1943],s[1942]} = (x[1942]+y[1942]+z[1942]);
assign {c[1944],s[1943]} = (x[1943]+y[1943]+z[1943]);
assign {c[1945],s[1944]} = (x[1944]+y[1944]+z[1944]);
assign {c[1946],s[1945]} = (x[1945]+y[1945]+z[1945]);
assign {c[1947],s[1946]} = (x[1946]+y[1946]+z[1946]);
assign {c[1948],s[1947]} = (x[1947]+y[1947]+z[1947]);
assign {c[1949],s[1948]} = (x[1948]+y[1948]+z[1948]);
assign {c[1950],s[1949]} = (x[1949]+y[1949]+z[1949]);
assign {c[1951],s[1950]} = (x[1950]+y[1950]+z[1950]);
assign {c[1952],s[1951]} = (x[1951]+y[1951]+z[1951]);
assign {c[1953],s[1952]} = (x[1952]+y[1952]+z[1952]);
assign {c[1954],s[1953]} = (x[1953]+y[1953]+z[1953]);
assign {c[1955],s[1954]} = (x[1954]+y[1954]+z[1954]);
assign {c[1956],s[1955]} = (x[1955]+y[1955]+z[1955]);
assign {c[1957],s[1956]} = (x[1956]+y[1956]+z[1956]);
assign {c[1958],s[1957]} = (x[1957]+y[1957]+z[1957]);
assign {c[1959],s[1958]} = (x[1958]+y[1958]+z[1958]);
assign {c[1960],s[1959]} = (x[1959]+y[1959]+z[1959]);
assign {c[1961],s[1960]} = (x[1960]+y[1960]+z[1960]);
assign {c[1962],s[1961]} = (x[1961]+y[1961]+z[1961]);
assign {c[1963],s[1962]} = (x[1962]+y[1962]+z[1962]);
assign {c[1964],s[1963]} = (x[1963]+y[1963]+z[1963]);
assign {c[1965],s[1964]} = (x[1964]+y[1964]+z[1964]);
assign {c[1966],s[1965]} = (x[1965]+y[1965]+z[1965]);
assign {c[1967],s[1966]} = (x[1966]+y[1966]+z[1966]);
assign {c[1968],s[1967]} = (x[1967]+y[1967]+z[1967]);
assign {c[1969],s[1968]} = (x[1968]+y[1968]+z[1968]);
assign {c[1970],s[1969]} = (x[1969]+y[1969]+z[1969]);
assign {c[1971],s[1970]} = (x[1970]+y[1970]+z[1970]);
assign {c[1972],s[1971]} = (x[1971]+y[1971]+z[1971]);
assign {c[1973],s[1972]} = (x[1972]+y[1972]+z[1972]);
assign {c[1974],s[1973]} = (x[1973]+y[1973]+z[1973]);
assign {c[1975],s[1974]} = (x[1974]+y[1974]+z[1974]);
assign {c[1976],s[1975]} = (x[1975]+y[1975]+z[1975]);
assign {c[1977],s[1976]} = (x[1976]+y[1976]+z[1976]);
assign {c[1978],s[1977]} = (x[1977]+y[1977]+z[1977]);
assign {c[1979],s[1978]} = (x[1978]+y[1978]+z[1978]);
assign {c[1980],s[1979]} = (x[1979]+y[1979]+z[1979]);
assign {c[1981],s[1980]} = (x[1980]+y[1980]+z[1980]);
assign {c[1982],s[1981]} = (x[1981]+y[1981]+z[1981]);
assign {c[1983],s[1982]} = (x[1982]+y[1982]+z[1982]);
assign {c[1984],s[1983]} = (x[1983]+y[1983]+z[1983]);
assign {c[1985],s[1984]} = (x[1984]+y[1984]+z[1984]);
assign {c[1986],s[1985]} = (x[1985]+y[1985]+z[1985]);
assign {c[1987],s[1986]} = (x[1986]+y[1986]+z[1986]);
assign {c[1988],s[1987]} = (x[1987]+y[1987]+z[1987]);
assign {c[1989],s[1988]} = (x[1988]+y[1988]+z[1988]);
assign {c[1990],s[1989]} = (x[1989]+y[1989]+z[1989]);
assign {c[1991],s[1990]} = (x[1990]+y[1990]+z[1990]);
assign {c[1992],s[1991]} = (x[1991]+y[1991]+z[1991]);
assign {c[1993],s[1992]} = (x[1992]+y[1992]+z[1992]);
assign {c[1994],s[1993]} = (x[1993]+y[1993]+z[1993]);
assign {c[1995],s[1994]} = (x[1994]+y[1994]+z[1994]);
assign {c[1996],s[1995]} = (x[1995]+y[1995]+z[1995]);
assign {c[1997],s[1996]} = (x[1996]+y[1996]+z[1996]);
assign {c[1998],s[1997]} = (x[1997]+y[1997]+z[1997]);
assign {c[1999],s[1998]} = (x[1998]+y[1998]+z[1998]);
assign {c[2000],s[1999]} = (x[1999]+y[1999]+z[1999]);
assign {c[2001],s[2000]} = (x[2000]+y[2000]+z[2000]);
assign {c[2002],s[2001]} = (x[2001]+y[2001]+z[2001]);
assign {c[2003],s[2002]} = (x[2002]+y[2002]+z[2002]);
assign {c[2004],s[2003]} = (x[2003]+y[2003]+z[2003]);
assign {c[2005],s[2004]} = (x[2004]+y[2004]+z[2004]);
assign {c[2006],s[2005]} = (x[2005]+y[2005]+z[2005]);
assign {c[2007],s[2006]} = (x[2006]+y[2006]+z[2006]);
assign {c[2008],s[2007]} = (x[2007]+y[2007]+z[2007]);
assign {c[2009],s[2008]} = (x[2008]+y[2008]+z[2008]);
assign {c[2010],s[2009]} = (x[2009]+y[2009]+z[2009]);
assign {c[2011],s[2010]} = (x[2010]+y[2010]+z[2010]);
assign {c[2012],s[2011]} = (x[2011]+y[2011]+z[2011]);
assign {c[2013],s[2012]} = (x[2012]+y[2012]+z[2012]);
assign {c[2014],s[2013]} = (x[2013]+y[2013]+z[2013]);
assign {c[2015],s[2014]} = (x[2014]+y[2014]+z[2014]);
assign {c[2016],s[2015]} = (x[2015]+y[2015]+z[2015]);
assign {c[2017],s[2016]} = (x[2016]+y[2016]+z[2016]);
assign {c[2018],s[2017]} = (x[2017]+y[2017]+z[2017]);
assign {c[2019],s[2018]} = (x[2018]+y[2018]+z[2018]);
assign {c[2020],s[2019]} = (x[2019]+y[2019]+z[2019]);
assign {c[2021],s[2020]} = (x[2020]+y[2020]+z[2020]);
assign {c[2022],s[2021]} = (x[2021]+y[2021]+z[2021]);
assign {c[2023],s[2022]} = (x[2022]+y[2022]+z[2022]);
assign {c[2024],s[2023]} = (x[2023]+y[2023]+z[2023]);
assign {c[2025],s[2024]} = (x[2024]+y[2024]+z[2024]);
assign {c[2026],s[2025]} = (x[2025]+y[2025]+z[2025]);
assign {c[2027],s[2026]} = (x[2026]+y[2026]+z[2026]);
assign {c[2028],s[2027]} = (x[2027]+y[2027]+z[2027]);
assign {c[2029],s[2028]} = (x[2028]+y[2028]+z[2028]);
assign {c[2030],s[2029]} = (x[2029]+y[2029]+z[2029]);
assign {c[2031],s[2030]} = (x[2030]+y[2030]+z[2030]);
assign {c[2032],s[2031]} = (x[2031]+y[2031]+z[2031]);
assign {c[2033],s[2032]} = (x[2032]+y[2032]+z[2032]);
assign {c[2034],s[2033]} = (x[2033]+y[2033]+z[2033]);
assign {c[2035],s[2034]} = (x[2034]+y[2034]+z[2034]);
assign {c[2036],s[2035]} = (x[2035]+y[2035]+z[2035]);
assign {c[2037],s[2036]} = (x[2036]+y[2036]+z[2036]);
assign {c[2038],s[2037]} = (x[2037]+y[2037]+z[2037]);
assign {c[2039],s[2038]} = (x[2038]+y[2038]+z[2038]);
assign {c[2040],s[2039]} = (x[2039]+y[2039]+z[2039]);
assign {c[2041],s[2040]} = (x[2040]+y[2040]+z[2040]);
assign {c[2042],s[2041]} = (x[2041]+y[2041]+z[2041]);
assign {c[2043],s[2042]} = (x[2042]+y[2042]+z[2042]);
assign {c[2044],s[2043]} = (x[2043]+y[2043]+z[2043]);
assign {c[2045],s[2044]} = (x[2044]+y[2044]+z[2044]);
assign {c[2046],s[2045]} = (x[2045]+y[2045]+z[2045]);
assign {c[2047],s[2046]} = (x[2046]+y[2046]+z[2046]);
assign {c[2048],s[2047]} = (x[2047]+y[2047]+z[2047]);
assign {c[2049],s[2048]} = (x[2048]+y[2048]+z[2048]);
assign {c[2050],s[2049]} = (x[2049]+y[2049]+z[2049]);
assign {c[2051],s[2050]} = (x[2050]+y[2050]+z[2050]);
assign {c[2052],s[2051]} = (x[2051]+y[2051]+z[2051]);
assign {c[2053],s[2052]} = (x[2052]+y[2052]+z[2052]);
assign {c[2054],s[2053]} = (x[2053]+y[2053]+z[2053]);
assign {c[2055],s[2054]} = (x[2054]+y[2054]+z[2054]);
assign {c[2056],s[2055]} = (x[2055]+y[2055]+z[2055]);
assign {c[2057],s[2056]} = (x[2056]+y[2056]+z[2056]);
assign {c[2058],s[2057]} = (x[2057]+y[2057]+z[2057]);
assign {c[2059],s[2058]} = (x[2058]+y[2058]+z[2058]);
assign {c[2060],s[2059]} = (x[2059]+y[2059]+z[2059]);
assign {c[2061],s[2060]} = (x[2060]+y[2060]+z[2060]);
assign {c[2062],s[2061]} = (x[2061]+y[2061]+z[2061]);
assign {c[2063],s[2062]} = (x[2062]+y[2062]+z[2062]);
assign {c[2064],s[2063]} = (x[2063]+y[2063]+z[2063]);
assign {c[2065],s[2064]} = (x[2064]+y[2064]+z[2064]);
assign {c[2066],s[2065]} = (x[2065]+y[2065]+z[2065]);
assign {c[2067],s[2066]} = (x[2066]+y[2066]+z[2066]);
assign {c[2068],s[2067]} = (x[2067]+y[2067]+z[2067]);
assign {c[2069],s[2068]} = (x[2068]+y[2068]+z[2068]);
assign {c[2070],s[2069]} = (x[2069]+y[2069]+z[2069]);
assign {c[2071],s[2070]} = (x[2070]+y[2070]+z[2070]);
assign {c[2072],s[2071]} = (x[2071]+y[2071]+z[2071]);
assign {c[2073],s[2072]} = (x[2072]+y[2072]+z[2072]);
assign {c[2074],s[2073]} = (x[2073]+y[2073]+z[2073]);
assign {c[2075],s[2074]} = (x[2074]+y[2074]+z[2074]);
assign {c[2076],s[2075]} = (x[2075]+y[2075]+z[2075]);
assign {c[2077],s[2076]} = (x[2076]+y[2076]+z[2076]);
assign {c[2078],s[2077]} = (x[2077]+y[2077]+z[2077]);
assign {c[2079],s[2078]} = (x[2078]+y[2078]+z[2078]);
assign {c[2080],s[2079]} = (x[2079]+y[2079]+z[2079]);
assign {c[2081],s[2080]} = (x[2080]+y[2080]+z[2080]);
assign {c[2082],s[2081]} = (x[2081]+y[2081]+z[2081]);
assign {c[2083],s[2082]} = (x[2082]+y[2082]+z[2082]);
assign {c[2084],s[2083]} = (x[2083]+y[2083]+z[2083]);
assign {c[2085],s[2084]} = (x[2084]+y[2084]+z[2084]);
assign {c[2086],s[2085]} = (x[2085]+y[2085]+z[2085]);
assign {c[2087],s[2086]} = (x[2086]+y[2086]+z[2086]);
assign {c[2088],s[2087]} = (x[2087]+y[2087]+z[2087]);
assign {c[2089],s[2088]} = (x[2088]+y[2088]+z[2088]);
assign {c[2090],s[2089]} = (x[2089]+y[2089]+z[2089]);
assign {c[2091],s[2090]} = (x[2090]+y[2090]+z[2090]);
assign {c[2092],s[2091]} = (x[2091]+y[2091]+z[2091]);
assign {c[2093],s[2092]} = (x[2092]+y[2092]+z[2092]);
assign {c[2094],s[2093]} = (x[2093]+y[2093]+z[2093]);
assign {c[2095],s[2094]} = (x[2094]+y[2094]+z[2094]);
assign {c[2096],s[2095]} = (x[2095]+y[2095]+z[2095]);
assign {c[2097],s[2096]} = (x[2096]+y[2096]+z[2096]);
assign {c[2098],s[2097]} = (x[2097]+y[2097]+z[2097]);
assign {c[2099],s[2098]} = (x[2098]+y[2098]+z[2098]);
assign {c[2100],s[2099]} = (x[2099]+y[2099]+z[2099]);
assign {c[2101],s[2100]} = (x[2100]+y[2100]+z[2100]);
assign {c[2102],s[2101]} = (x[2101]+y[2101]+z[2101]);
assign {c[2103],s[2102]} = (x[2102]+y[2102]+z[2102]);
assign {c[2104],s[2103]} = (x[2103]+y[2103]+z[2103]);
assign {c[2105],s[2104]} = (x[2104]+y[2104]+z[2104]);
assign {c[2106],s[2105]} = (x[2105]+y[2105]+z[2105]);
assign {c[2107],s[2106]} = (x[2106]+y[2106]+z[2106]);
assign {c[2108],s[2107]} = (x[2107]+y[2107]+z[2107]);
assign {c[2109],s[2108]} = (x[2108]+y[2108]+z[2108]);
assign {c[2110],s[2109]} = (x[2109]+y[2109]+z[2109]);
assign {c[2111],s[2110]} = (x[2110]+y[2110]+z[2110]);
assign {c[2112],s[2111]} = (x[2111]+y[2111]+z[2111]);
assign {c[2113],s[2112]} = (x[2112]+y[2112]+z[2112]);
assign {c[2114],s[2113]} = (x[2113]+y[2113]+z[2113]);
assign {c[2115],s[2114]} = (x[2114]+y[2114]+z[2114]);
assign {c[2116],s[2115]} = (x[2115]+y[2115]+z[2115]);
assign {c[2117],s[2116]} = (x[2116]+y[2116]+z[2116]);
assign {c[2118],s[2117]} = (x[2117]+y[2117]+z[2117]);
assign {c[2119],s[2118]} = (x[2118]+y[2118]+z[2118]);
assign {c[2120],s[2119]} = (x[2119]+y[2119]+z[2119]);
assign {c[2121],s[2120]} = (x[2120]+y[2120]+z[2120]);
assign {c[2122],s[2121]} = (x[2121]+y[2121]+z[2121]);
assign {c[2123],s[2122]} = (x[2122]+y[2122]+z[2122]);
assign {c[2124],s[2123]} = (x[2123]+y[2123]+z[2123]);
assign {c[2125],s[2124]} = (x[2124]+y[2124]+z[2124]);
assign {c[2126],s[2125]} = (x[2125]+y[2125]+z[2125]);
assign {c[2127],s[2126]} = (x[2126]+y[2126]+z[2126]);
assign {c[2128],s[2127]} = (x[2127]+y[2127]+z[2127]);
assign {c[2129],s[2128]} = (x[2128]+y[2128]+z[2128]);
assign {c[2130],s[2129]} = (x[2129]+y[2129]+z[2129]);
assign {c[2131],s[2130]} = (x[2130]+y[2130]+z[2130]);
assign {c[2132],s[2131]} = (x[2131]+y[2131]+z[2131]);
assign {c[2133],s[2132]} = (x[2132]+y[2132]+z[2132]);
assign {c[2134],s[2133]} = (x[2133]+y[2133]+z[2133]);
assign {c[2135],s[2134]} = (x[2134]+y[2134]+z[2134]);
assign {c[2136],s[2135]} = (x[2135]+y[2135]+z[2135]);
assign {c[2137],s[2136]} = (x[2136]+y[2136]+z[2136]);
assign {c[2138],s[2137]} = (x[2137]+y[2137]+z[2137]);
assign {c[2139],s[2138]} = (x[2138]+y[2138]+z[2138]);
assign {c[2140],s[2139]} = (x[2139]+y[2139]+z[2139]);
assign {c[2141],s[2140]} = (x[2140]+y[2140]+z[2140]);
assign {c[2142],s[2141]} = (x[2141]+y[2141]+z[2141]);
assign {c[2143],s[2142]} = (x[2142]+y[2142]+z[2142]);
assign {c[2144],s[2143]} = (x[2143]+y[2143]+z[2143]);
assign {c[2145],s[2144]} = (x[2144]+y[2144]+z[2144]);
assign {c[2146],s[2145]} = (x[2145]+y[2145]+z[2145]);
assign {c[2147],s[2146]} = (x[2146]+y[2146]+z[2146]);
assign {c[2148],s[2147]} = (x[2147]+y[2147]+z[2147]);
assign {c[2149],s[2148]} = (x[2148]+y[2148]+z[2148]);
assign {c[2150],s[2149]} = (x[2149]+y[2149]+z[2149]);
assign {c[2151],s[2150]} = (x[2150]+y[2150]+z[2150]);
assign {c[2152],s[2151]} = (x[2151]+y[2151]+z[2151]);
assign {c[2153],s[2152]} = (x[2152]+y[2152]+z[2152]);
assign {c[2154],s[2153]} = (x[2153]+y[2153]+z[2153]);
assign {c[2155],s[2154]} = (x[2154]+y[2154]+z[2154]);
assign {c[2156],s[2155]} = (x[2155]+y[2155]+z[2155]);
assign {c[2157],s[2156]} = (x[2156]+y[2156]+z[2156]);
assign {c[2158],s[2157]} = (x[2157]+y[2157]+z[2157]);
assign {c[2159],s[2158]} = (x[2158]+y[2158]+z[2158]);
assign {c[2160],s[2159]} = (x[2159]+y[2159]+z[2159]);
assign {c[2161],s[2160]} = (x[2160]+y[2160]+z[2160]);
assign {c[2162],s[2161]} = (x[2161]+y[2161]+z[2161]);
assign {c[2163],s[2162]} = (x[2162]+y[2162]+z[2162]);
assign {c[2164],s[2163]} = (x[2163]+y[2163]+z[2163]);
assign {c[2165],s[2164]} = (x[2164]+y[2164]+z[2164]);
assign {c[2166],s[2165]} = (x[2165]+y[2165]+z[2165]);
assign {c[2167],s[2166]} = (x[2166]+y[2166]+z[2166]);
assign {c[2168],s[2167]} = (x[2167]+y[2167]+z[2167]);
assign {c[2169],s[2168]} = (x[2168]+y[2168]+z[2168]);
assign {c[2170],s[2169]} = (x[2169]+y[2169]+z[2169]);
assign {c[2171],s[2170]} = (x[2170]+y[2170]+z[2170]);
assign {c[2172],s[2171]} = (x[2171]+y[2171]+z[2171]);
assign {c[2173],s[2172]} = (x[2172]+y[2172]+z[2172]);
assign {c[2174],s[2173]} = (x[2173]+y[2173]+z[2173]);
assign {c[2175],s[2174]} = (x[2174]+y[2174]+z[2174]);
assign {c[2176],s[2175]} = (x[2175]+y[2175]+z[2175]);
assign {c[2177],s[2176]} = (x[2176]+y[2176]+z[2176]);
assign {c[2178],s[2177]} = (x[2177]+y[2177]+z[2177]);
assign {c[2179],s[2178]} = (x[2178]+y[2178]+z[2178]);
assign {c[2180],s[2179]} = (x[2179]+y[2179]+z[2179]);
assign {c[2181],s[2180]} = (x[2180]+y[2180]+z[2180]);
assign {c[2182],s[2181]} = (x[2181]+y[2181]+z[2181]);
assign {c[2183],s[2182]} = (x[2182]+y[2182]+z[2182]);
assign {c[2184],s[2183]} = (x[2183]+y[2183]+z[2183]);
assign {c[2185],s[2184]} = (x[2184]+y[2184]+z[2184]);
assign {c[2186],s[2185]} = (x[2185]+y[2185]+z[2185]);
assign {c[2187],s[2186]} = (x[2186]+y[2186]+z[2186]);
assign {c[2188],s[2187]} = (x[2187]+y[2187]+z[2187]);
assign {c[2189],s[2188]} = (x[2188]+y[2188]+z[2188]);
assign {c[2190],s[2189]} = (x[2189]+y[2189]+z[2189]);
assign {c[2191],s[2190]} = (x[2190]+y[2190]+z[2190]);
assign {c[2192],s[2191]} = (x[2191]+y[2191]+z[2191]);
assign {c[2193],s[2192]} = (x[2192]+y[2192]+z[2192]);
assign {c[2194],s[2193]} = (x[2193]+y[2193]+z[2193]);
assign {c[2195],s[2194]} = (x[2194]+y[2194]+z[2194]);
assign {c[2196],s[2195]} = (x[2195]+y[2195]+z[2195]);
assign {c[2197],s[2196]} = (x[2196]+y[2196]+z[2196]);
assign {c[2198],s[2197]} = (x[2197]+y[2197]+z[2197]);
assign {c[2199],s[2198]} = (x[2198]+y[2198]+z[2198]);
assign {c[2200],s[2199]} = (x[2199]+y[2199]+z[2199]);
assign {c[2201],s[2200]} = (x[2200]+y[2200]+z[2200]);
assign {c[2202],s[2201]} = (x[2201]+y[2201]+z[2201]);
assign {c[2203],s[2202]} = (x[2202]+y[2202]+z[2202]);
assign {c[2204],s[2203]} = (x[2203]+y[2203]+z[2203]);
assign {c[2205],s[2204]} = (x[2204]+y[2204]+z[2204]);
assign {c[2206],s[2205]} = (x[2205]+y[2205]+z[2205]);
assign {c[2207],s[2206]} = (x[2206]+y[2206]+z[2206]);
assign {c[2208],s[2207]} = (x[2207]+y[2207]+z[2207]);
assign {c[2209],s[2208]} = (x[2208]+y[2208]+z[2208]);
assign {c[2210],s[2209]} = (x[2209]+y[2209]+z[2209]);
assign {c[2211],s[2210]} = (x[2210]+y[2210]+z[2210]);
assign {c[2212],s[2211]} = (x[2211]+y[2211]+z[2211]);
assign {c[2213],s[2212]} = (x[2212]+y[2212]+z[2212]);
assign {c[2214],s[2213]} = (x[2213]+y[2213]+z[2213]);
assign {c[2215],s[2214]} = (x[2214]+y[2214]+z[2214]);
assign {c[2216],s[2215]} = (x[2215]+y[2215]+z[2215]);
assign {c[2217],s[2216]} = (x[2216]+y[2216]+z[2216]);
assign {c[2218],s[2217]} = (x[2217]+y[2217]+z[2217]);
assign {c[2219],s[2218]} = (x[2218]+y[2218]+z[2218]);
assign {c[2220],s[2219]} = (x[2219]+y[2219]+z[2219]);
assign {c[2221],s[2220]} = (x[2220]+y[2220]+z[2220]);
assign {c[2222],s[2221]} = (x[2221]+y[2221]+z[2221]);
assign {c[2223],s[2222]} = (x[2222]+y[2222]+z[2222]);
assign {c[2224],s[2223]} = (x[2223]+y[2223]+z[2223]);
assign {c[2225],s[2224]} = (x[2224]+y[2224]+z[2224]);
assign {c[2226],s[2225]} = (x[2225]+y[2225]+z[2225]);
assign {c[2227],s[2226]} = (x[2226]+y[2226]+z[2226]);
assign {c[2228],s[2227]} = (x[2227]+y[2227]+z[2227]);
assign {c[2229],s[2228]} = (x[2228]+y[2228]+z[2228]);
assign {c[2230],s[2229]} = (x[2229]+y[2229]+z[2229]);
assign {c[2231],s[2230]} = (x[2230]+y[2230]+z[2230]);
assign {c[2232],s[2231]} = (x[2231]+y[2231]+z[2231]);
assign {c[2233],s[2232]} = (x[2232]+y[2232]+z[2232]);
assign {c[2234],s[2233]} = (x[2233]+y[2233]+z[2233]);
assign {c[2235],s[2234]} = (x[2234]+y[2234]+z[2234]);
assign {c[2236],s[2235]} = (x[2235]+y[2235]+z[2235]);
assign {c[2237],s[2236]} = (x[2236]+y[2236]+z[2236]);
assign {c[2238],s[2237]} = (x[2237]+y[2237]+z[2237]);
assign {c[2239],s[2238]} = (x[2238]+y[2238]+z[2238]);
assign {c[2240],s[2239]} = (x[2239]+y[2239]+z[2239]);
assign {c[2241],s[2240]} = (x[2240]+y[2240]+z[2240]);
assign {c[2242],s[2241]} = (x[2241]+y[2241]+z[2241]);
assign {c[2243],s[2242]} = (x[2242]+y[2242]+z[2242]);
assign {c[2244],s[2243]} = (x[2243]+y[2243]+z[2243]);
assign {c[2245],s[2244]} = (x[2244]+y[2244]+z[2244]);
assign {c[2246],s[2245]} = (x[2245]+y[2245]+z[2245]);
assign {c[2247],s[2246]} = (x[2246]+y[2246]+z[2246]);
assign {c[2248],s[2247]} = (x[2247]+y[2247]+z[2247]);
assign {c[2249],s[2248]} = (x[2248]+y[2248]+z[2248]);
assign {c[2250],s[2249]} = (x[2249]+y[2249]+z[2249]);
assign {c[2251],s[2250]} = (x[2250]+y[2250]+z[2250]);
assign {c[2252],s[2251]} = (x[2251]+y[2251]+z[2251]);
assign {c[2253],s[2252]} = (x[2252]+y[2252]+z[2252]);
assign {c[2254],s[2253]} = (x[2253]+y[2253]+z[2253]);
assign {c[2255],s[2254]} = (x[2254]+y[2254]+z[2254]);
assign {c[2256],s[2255]} = (x[2255]+y[2255]+z[2255]);
assign {c[2257],s[2256]} = (x[2256]+y[2256]+z[2256]);
assign {c[2258],s[2257]} = (x[2257]+y[2257]+z[2257]);
assign {c[2259],s[2258]} = (x[2258]+y[2258]+z[2258]);
assign {c[2260],s[2259]} = (x[2259]+y[2259]+z[2259]);
assign {c[2261],s[2260]} = (x[2260]+y[2260]+z[2260]);
assign {c[2262],s[2261]} = (x[2261]+y[2261]+z[2261]);
assign {c[2263],s[2262]} = (x[2262]+y[2262]+z[2262]);
assign {c[2264],s[2263]} = (x[2263]+y[2263]+z[2263]);
assign {c[2265],s[2264]} = (x[2264]+y[2264]+z[2264]);
assign {c[2266],s[2265]} = (x[2265]+y[2265]+z[2265]);
assign {c[2267],s[2266]} = (x[2266]+y[2266]+z[2266]);
assign {c[2268],s[2267]} = (x[2267]+y[2267]+z[2267]);
assign {c[2269],s[2268]} = (x[2268]+y[2268]+z[2268]);
assign {c[2270],s[2269]} = (x[2269]+y[2269]+z[2269]);
assign {c[2271],s[2270]} = (x[2270]+y[2270]+z[2270]);
assign {c[2272],s[2271]} = (x[2271]+y[2271]+z[2271]);
assign {c[2273],s[2272]} = (x[2272]+y[2272]+z[2272]);
assign {c[2274],s[2273]} = (x[2273]+y[2273]+z[2273]);
assign {c[2275],s[2274]} = (x[2274]+y[2274]+z[2274]);
assign {c[2276],s[2275]} = (x[2275]+y[2275]+z[2275]);
assign {c[2277],s[2276]} = (x[2276]+y[2276]+z[2276]);
assign {c[2278],s[2277]} = (x[2277]+y[2277]+z[2277]);
assign {c[2279],s[2278]} = (x[2278]+y[2278]+z[2278]);
assign {c[2280],s[2279]} = (x[2279]+y[2279]+z[2279]);
assign {c[2281],s[2280]} = (x[2280]+y[2280]+z[2280]);
assign {c[2282],s[2281]} = (x[2281]+y[2281]+z[2281]);
assign {c[2283],s[2282]} = (x[2282]+y[2282]+z[2282]);
assign {c[2284],s[2283]} = (x[2283]+y[2283]+z[2283]);
assign {c[2285],s[2284]} = (x[2284]+y[2284]+z[2284]);
assign {c[2286],s[2285]} = (x[2285]+y[2285]+z[2285]);
assign {c[2287],s[2286]} = (x[2286]+y[2286]+z[2286]);
assign {c[2288],s[2287]} = (x[2287]+y[2287]+z[2287]);
assign {c[2289],s[2288]} = (x[2288]+y[2288]+z[2288]);
assign {c[2290],s[2289]} = (x[2289]+y[2289]+z[2289]);
assign {c[2291],s[2290]} = (x[2290]+y[2290]+z[2290]);
assign {c[2292],s[2291]} = (x[2291]+y[2291]+z[2291]);
assign {c[2293],s[2292]} = (x[2292]+y[2292]+z[2292]);
assign {c[2294],s[2293]} = (x[2293]+y[2293]+z[2293]);
assign {c[2295],s[2294]} = (x[2294]+y[2294]+z[2294]);
assign {c[2296],s[2295]} = (x[2295]+y[2295]+z[2295]);
assign {c[2297],s[2296]} = (x[2296]+y[2296]+z[2296]);
assign {c[2298],s[2297]} = (x[2297]+y[2297]+z[2297]);
assign {c[2299],s[2298]} = (x[2298]+y[2298]+z[2298]);
assign {c[2300],s[2299]} = (x[2299]+y[2299]+z[2299]);
assign {c[2301],s[2300]} = (x[2300]+y[2300]+z[2300]);
assign {c[2302],s[2301]} = (x[2301]+y[2301]+z[2301]);
assign {c[2303],s[2302]} = (x[2302]+y[2302]+z[2302]);
assign {c[2304],s[2303]} = (x[2303]+y[2303]+z[2303]);
assign {c[2305],s[2304]} = (x[2304]+y[2304]+z[2304]);
assign {c[2306],s[2305]} = (x[2305]+y[2305]+z[2305]);
assign {c[2307],s[2306]} = (x[2306]+y[2306]+z[2306]);
assign {c[2308],s[2307]} = (x[2307]+y[2307]+z[2307]);
assign {c[2309],s[2308]} = (x[2308]+y[2308]+z[2308]);
assign {c[2310],s[2309]} = (x[2309]+y[2309]+z[2309]);
assign {c[2311],s[2310]} = (x[2310]+y[2310]+z[2310]);
assign {c[2312],s[2311]} = (x[2311]+y[2311]+z[2311]);
assign {c[2313],s[2312]} = (x[2312]+y[2312]+z[2312]);
assign {c[2314],s[2313]} = (x[2313]+y[2313]+z[2313]);
assign {c[2315],s[2314]} = (x[2314]+y[2314]+z[2314]);
assign {c[2316],s[2315]} = (x[2315]+y[2315]+z[2315]);
assign {c[2317],s[2316]} = (x[2316]+y[2316]+z[2316]);
assign {c[2318],s[2317]} = (x[2317]+y[2317]+z[2317]);
assign {c[2319],s[2318]} = (x[2318]+y[2318]+z[2318]);
assign {c[2320],s[2319]} = (x[2319]+y[2319]+z[2319]);
assign {c[2321],s[2320]} = (x[2320]+y[2320]+z[2320]);
assign {c[2322],s[2321]} = (x[2321]+y[2321]+z[2321]);
assign {c[2323],s[2322]} = (x[2322]+y[2322]+z[2322]);
assign {c[2324],s[2323]} = (x[2323]+y[2323]+z[2323]);
assign {c[2325],s[2324]} = (x[2324]+y[2324]+z[2324]);
assign {c[2326],s[2325]} = (x[2325]+y[2325]+z[2325]);
assign {c[2327],s[2326]} = (x[2326]+y[2326]+z[2326]);
assign {c[2328],s[2327]} = (x[2327]+y[2327]+z[2327]);
assign {c[2329],s[2328]} = (x[2328]+y[2328]+z[2328]);
assign {c[2330],s[2329]} = (x[2329]+y[2329]+z[2329]);
assign {c[2331],s[2330]} = (x[2330]+y[2330]+z[2330]);
assign {c[2332],s[2331]} = (x[2331]+y[2331]+z[2331]);
assign {c[2333],s[2332]} = (x[2332]+y[2332]+z[2332]);
assign {c[2334],s[2333]} = (x[2333]+y[2333]+z[2333]);
assign {c[2335],s[2334]} = (x[2334]+y[2334]+z[2334]);
assign {c[2336],s[2335]} = (x[2335]+y[2335]+z[2335]);
assign {c[2337],s[2336]} = (x[2336]+y[2336]+z[2336]);
assign {c[2338],s[2337]} = (x[2337]+y[2337]+z[2337]);
assign {c[2339],s[2338]} = (x[2338]+y[2338]+z[2338]);
assign {c[2340],s[2339]} = (x[2339]+y[2339]+z[2339]);
assign {c[2341],s[2340]} = (x[2340]+y[2340]+z[2340]);
assign {c[2342],s[2341]} = (x[2341]+y[2341]+z[2341]);
assign {c[2343],s[2342]} = (x[2342]+y[2342]+z[2342]);
assign {c[2344],s[2343]} = (x[2343]+y[2343]+z[2343]);
assign {c[2345],s[2344]} = (x[2344]+y[2344]+z[2344]);
assign {c[2346],s[2345]} = (x[2345]+y[2345]+z[2345]);
assign {c[2347],s[2346]} = (x[2346]+y[2346]+z[2346]);
assign {c[2348],s[2347]} = (x[2347]+y[2347]+z[2347]);
assign {c[2349],s[2348]} = (x[2348]+y[2348]+z[2348]);
assign {c[2350],s[2349]} = (x[2349]+y[2349]+z[2349]);
assign {c[2351],s[2350]} = (x[2350]+y[2350]+z[2350]);
assign {c[2352],s[2351]} = (x[2351]+y[2351]+z[2351]);
assign {c[2353],s[2352]} = (x[2352]+y[2352]+z[2352]);
assign {c[2354],s[2353]} = (x[2353]+y[2353]+z[2353]);
assign {c[2355],s[2354]} = (x[2354]+y[2354]+z[2354]);
assign {c[2356],s[2355]} = (x[2355]+y[2355]+z[2355]);
assign {c[2357],s[2356]} = (x[2356]+y[2356]+z[2356]);
assign {c[2358],s[2357]} = (x[2357]+y[2357]+z[2357]);
assign {c[2359],s[2358]} = (x[2358]+y[2358]+z[2358]);
assign {c[2360],s[2359]} = (x[2359]+y[2359]+z[2359]);
assign {c[2361],s[2360]} = (x[2360]+y[2360]+z[2360]);
assign {c[2362],s[2361]} = (x[2361]+y[2361]+z[2361]);
assign {c[2363],s[2362]} = (x[2362]+y[2362]+z[2362]);
assign {c[2364],s[2363]} = (x[2363]+y[2363]+z[2363]);
assign {c[2365],s[2364]} = (x[2364]+y[2364]+z[2364]);
assign {c[2366],s[2365]} = (x[2365]+y[2365]+z[2365]);
assign {c[2367],s[2366]} = (x[2366]+y[2366]+z[2366]);
assign {c[2368],s[2367]} = (x[2367]+y[2367]+z[2367]);
assign {c[2369],s[2368]} = (x[2368]+y[2368]+z[2368]);
assign {c[2370],s[2369]} = (x[2369]+y[2369]+z[2369]);
assign {c[2371],s[2370]} = (x[2370]+y[2370]+z[2370]);
assign {c[2372],s[2371]} = (x[2371]+y[2371]+z[2371]);
assign {c[2373],s[2372]} = (x[2372]+y[2372]+z[2372]);
assign {c[2374],s[2373]} = (x[2373]+y[2373]+z[2373]);
assign {c[2375],s[2374]} = (x[2374]+y[2374]+z[2374]);
assign {c[2376],s[2375]} = (x[2375]+y[2375]+z[2375]);
assign {c[2377],s[2376]} = (x[2376]+y[2376]+z[2376]);
assign {c[2378],s[2377]} = (x[2377]+y[2377]+z[2377]);
assign {c[2379],s[2378]} = (x[2378]+y[2378]+z[2378]);
assign {c[2380],s[2379]} = (x[2379]+y[2379]+z[2379]);
assign {c[2381],s[2380]} = (x[2380]+y[2380]+z[2380]);
assign {c[2382],s[2381]} = (x[2381]+y[2381]+z[2381]);
assign {c[2383],s[2382]} = (x[2382]+y[2382]+z[2382]);
assign {c[2384],s[2383]} = (x[2383]+y[2383]+z[2383]);
assign {c[2385],s[2384]} = (x[2384]+y[2384]+z[2384]);
assign {c[2386],s[2385]} = (x[2385]+y[2385]+z[2385]);
assign {c[2387],s[2386]} = (x[2386]+y[2386]+z[2386]);
assign {c[2388],s[2387]} = (x[2387]+y[2387]+z[2387]);
assign {c[2389],s[2388]} = (x[2388]+y[2388]+z[2388]);
assign {c[2390],s[2389]} = (x[2389]+y[2389]+z[2389]);
assign {c[2391],s[2390]} = (x[2390]+y[2390]+z[2390]);
assign {c[2392],s[2391]} = (x[2391]+y[2391]+z[2391]);
assign {c[2393],s[2392]} = (x[2392]+y[2392]+z[2392]);
assign {c[2394],s[2393]} = (x[2393]+y[2393]+z[2393]);
assign {c[2395],s[2394]} = (x[2394]+y[2394]+z[2394]);
assign {c[2396],s[2395]} = (x[2395]+y[2395]+z[2395]);
assign {c[2397],s[2396]} = (x[2396]+y[2396]+z[2396]);
assign {c[2398],s[2397]} = (x[2397]+y[2397]+z[2397]);
assign {c[2399],s[2398]} = (x[2398]+y[2398]+z[2398]);
assign {c[2400],s[2399]} = (x[2399]+y[2399]+z[2399]);
assign {c[2401],s[2400]} = (x[2400]+y[2400]+z[2400]);
assign {c[2402],s[2401]} = (x[2401]+y[2401]+z[2401]);
assign {c[2403],s[2402]} = (x[2402]+y[2402]+z[2402]);
assign {c[2404],s[2403]} = (x[2403]+y[2403]+z[2403]);
assign {c[2405],s[2404]} = (x[2404]+y[2404]+z[2404]);
assign {c[2406],s[2405]} = (x[2405]+y[2405]+z[2405]);
assign {c[2407],s[2406]} = (x[2406]+y[2406]+z[2406]);
assign {c[2408],s[2407]} = (x[2407]+y[2407]+z[2407]);
assign {c[2409],s[2408]} = (x[2408]+y[2408]+z[2408]);
assign {c[2410],s[2409]} = (x[2409]+y[2409]+z[2409]);
assign {c[2411],s[2410]} = (x[2410]+y[2410]+z[2410]);
assign {c[2412],s[2411]} = (x[2411]+y[2411]+z[2411]);
assign {c[2413],s[2412]} = (x[2412]+y[2412]+z[2412]);
assign {c[2414],s[2413]} = (x[2413]+y[2413]+z[2413]);
assign {c[2415],s[2414]} = (x[2414]+y[2414]+z[2414]);
assign {c[2416],s[2415]} = (x[2415]+y[2415]+z[2415]);
assign {c[2417],s[2416]} = (x[2416]+y[2416]+z[2416]);
assign {c[2418],s[2417]} = (x[2417]+y[2417]+z[2417]);
assign {c[2419],s[2418]} = (x[2418]+y[2418]+z[2418]);
assign {c[2420],s[2419]} = (x[2419]+y[2419]+z[2419]);
assign {c[2421],s[2420]} = (x[2420]+y[2420]+z[2420]);
assign {c[2422],s[2421]} = (x[2421]+y[2421]+z[2421]);
assign {c[2423],s[2422]} = (x[2422]+y[2422]+z[2422]);
assign {c[2424],s[2423]} = (x[2423]+y[2423]+z[2423]);
assign {c[2425],s[2424]} = (x[2424]+y[2424]+z[2424]);
assign {c[2426],s[2425]} = (x[2425]+y[2425]+z[2425]);
assign {c[2427],s[2426]} = (x[2426]+y[2426]+z[2426]);
assign {c[2428],s[2427]} = (x[2427]+y[2427]+z[2427]);
assign {c[2429],s[2428]} = (x[2428]+y[2428]+z[2428]);
assign {c[2430],s[2429]} = (x[2429]+y[2429]+z[2429]);
assign {c[2431],s[2430]} = (x[2430]+y[2430]+z[2430]);
assign {c[2432],s[2431]} = (x[2431]+y[2431]+z[2431]);
assign {c[2433],s[2432]} = (x[2432]+y[2432]+z[2432]);
assign {c[2434],s[2433]} = (x[2433]+y[2433]+z[2433]);
assign {c[2435],s[2434]} = (x[2434]+y[2434]+z[2434]);
assign {c[2436],s[2435]} = (x[2435]+y[2435]+z[2435]);
assign {c[2437],s[2436]} = (x[2436]+y[2436]+z[2436]);
assign {c[2438],s[2437]} = (x[2437]+y[2437]+z[2437]);
assign {c[2439],s[2438]} = (x[2438]+y[2438]+z[2438]);
assign {c[2440],s[2439]} = (x[2439]+y[2439]+z[2439]);
assign {c[2441],s[2440]} = (x[2440]+y[2440]+z[2440]);
assign {c[2442],s[2441]} = (x[2441]+y[2441]+z[2441]);
assign {c[2443],s[2442]} = (x[2442]+y[2442]+z[2442]);
assign {c[2444],s[2443]} = (x[2443]+y[2443]+z[2443]);
assign {c[2445],s[2444]} = (x[2444]+y[2444]+z[2444]);
assign {c[2446],s[2445]} = (x[2445]+y[2445]+z[2445]);
assign {c[2447],s[2446]} = (x[2446]+y[2446]+z[2446]);
assign {c[2448],s[2447]} = (x[2447]+y[2447]+z[2447]);
assign {c[2449],s[2448]} = (x[2448]+y[2448]+z[2448]);
assign {c[2450],s[2449]} = (x[2449]+y[2449]+z[2449]);
assign {c[2451],s[2450]} = (x[2450]+y[2450]+z[2450]);
assign {c[2452],s[2451]} = (x[2451]+y[2451]+z[2451]);
assign {c[2453],s[2452]} = (x[2452]+y[2452]+z[2452]);
assign {c[2454],s[2453]} = (x[2453]+y[2453]+z[2453]);
assign {c[2455],s[2454]} = (x[2454]+y[2454]+z[2454]);
assign {c[2456],s[2455]} = (x[2455]+y[2455]+z[2455]);
assign {c[2457],s[2456]} = (x[2456]+y[2456]+z[2456]);
assign {c[2458],s[2457]} = (x[2457]+y[2457]+z[2457]);
assign {c[2459],s[2458]} = (x[2458]+y[2458]+z[2458]);
assign {c[2460],s[2459]} = (x[2459]+y[2459]+z[2459]);
assign {c[2461],s[2460]} = (x[2460]+y[2460]+z[2460]);
assign {c[2462],s[2461]} = (x[2461]+y[2461]+z[2461]);
assign {c[2463],s[2462]} = (x[2462]+y[2462]+z[2462]);
assign {c[2464],s[2463]} = (x[2463]+y[2463]+z[2463]);
assign {c[2465],s[2464]} = (x[2464]+y[2464]+z[2464]);
assign {c[2466],s[2465]} = (x[2465]+y[2465]+z[2465]);
assign {c[2467],s[2466]} = (x[2466]+y[2466]+z[2466]);
assign {c[2468],s[2467]} = (x[2467]+y[2467]+z[2467]);
assign {c[2469],s[2468]} = (x[2468]+y[2468]+z[2468]);
assign {c[2470],s[2469]} = (x[2469]+y[2469]+z[2469]);
assign {c[2471],s[2470]} = (x[2470]+y[2470]+z[2470]);
assign {c[2472],s[2471]} = (x[2471]+y[2471]+z[2471]);
assign {c[2473],s[2472]} = (x[2472]+y[2472]+z[2472]);
assign {c[2474],s[2473]} = (x[2473]+y[2473]+z[2473]);
assign {c[2475],s[2474]} = (x[2474]+y[2474]+z[2474]);
assign {c[2476],s[2475]} = (x[2475]+y[2475]+z[2475]);
assign {c[2477],s[2476]} = (x[2476]+y[2476]+z[2476]);
assign {c[2478],s[2477]} = (x[2477]+y[2477]+z[2477]);
assign {c[2479],s[2478]} = (x[2478]+y[2478]+z[2478]);
assign {c[2480],s[2479]} = (x[2479]+y[2479]+z[2479]);
assign {c[2481],s[2480]} = (x[2480]+y[2480]+z[2480]);
assign {c[2482],s[2481]} = (x[2481]+y[2481]+z[2481]);
assign {c[2483],s[2482]} = (x[2482]+y[2482]+z[2482]);
assign {c[2484],s[2483]} = (x[2483]+y[2483]+z[2483]);
assign {c[2485],s[2484]} = (x[2484]+y[2484]+z[2484]);
assign {c[2486],s[2485]} = (x[2485]+y[2485]+z[2485]);
assign {c[2487],s[2486]} = (x[2486]+y[2486]+z[2486]);
assign {c[2488],s[2487]} = (x[2487]+y[2487]+z[2487]);
assign {c[2489],s[2488]} = (x[2488]+y[2488]+z[2488]);
assign {c[2490],s[2489]} = (x[2489]+y[2489]+z[2489]);
assign {c[2491],s[2490]} = (x[2490]+y[2490]+z[2490]);
assign {c[2492],s[2491]} = (x[2491]+y[2491]+z[2491]);
assign {c[2493],s[2492]} = (x[2492]+y[2492]+z[2492]);
assign {c[2494],s[2493]} = (x[2493]+y[2493]+z[2493]);
assign {c[2495],s[2494]} = (x[2494]+y[2494]+z[2494]);
assign {c[2496],s[2495]} = (x[2495]+y[2495]+z[2495]);
assign {c[2497],s[2496]} = (x[2496]+y[2496]+z[2496]);
assign {c[2498],s[2497]} = (x[2497]+y[2497]+z[2497]);
assign {c[2499],s[2498]} = (x[2498]+y[2498]+z[2498]);
assign {c[2500],s[2499]} = (x[2499]+y[2499]+z[2499]);
assign {c[2501],s[2500]} = (x[2500]+y[2500]+z[2500]);
assign {c[2502],s[2501]} = (x[2501]+y[2501]+z[2501]);
assign {c[2503],s[2502]} = (x[2502]+y[2502]+z[2502]);
assign {c[2504],s[2503]} = (x[2503]+y[2503]+z[2503]);
assign {c[2505],s[2504]} = (x[2504]+y[2504]+z[2504]);
assign {c[2506],s[2505]} = (x[2505]+y[2505]+z[2505]);
assign {c[2507],s[2506]} = (x[2506]+y[2506]+z[2506]);
assign {c[2508],s[2507]} = (x[2507]+y[2507]+z[2507]);
assign {c[2509],s[2508]} = (x[2508]+y[2508]+z[2508]);
assign {c[2510],s[2509]} = (x[2509]+y[2509]+z[2509]);
assign {c[2511],s[2510]} = (x[2510]+y[2510]+z[2510]);
assign {c[2512],s[2511]} = (x[2511]+y[2511]+z[2511]);
assign {c[2513],s[2512]} = (x[2512]+y[2512]+z[2512]);
assign {c[2514],s[2513]} = (x[2513]+y[2513]+z[2513]);
assign {c[2515],s[2514]} = (x[2514]+y[2514]+z[2514]);
assign {c[2516],s[2515]} = (x[2515]+y[2515]+z[2515]);
assign {c[2517],s[2516]} = (x[2516]+y[2516]+z[2516]);
assign {c[2518],s[2517]} = (x[2517]+y[2517]+z[2517]);
assign {c[2519],s[2518]} = (x[2518]+y[2518]+z[2518]);
assign {c[2520],s[2519]} = (x[2519]+y[2519]+z[2519]);
assign {c[2521],s[2520]} = (x[2520]+y[2520]+z[2520]);
assign {c[2522],s[2521]} = (x[2521]+y[2521]+z[2521]);
assign {c[2523],s[2522]} = (x[2522]+y[2522]+z[2522]);
assign {c[2524],s[2523]} = (x[2523]+y[2523]+z[2523]);
assign {c[2525],s[2524]} = (x[2524]+y[2524]+z[2524]);
assign {c[2526],s[2525]} = (x[2525]+y[2525]+z[2525]);
assign {c[2527],s[2526]} = (x[2526]+y[2526]+z[2526]);
assign {c[2528],s[2527]} = (x[2527]+y[2527]+z[2527]);
assign {c[2529],s[2528]} = (x[2528]+y[2528]+z[2528]);
assign {c[2530],s[2529]} = (x[2529]+y[2529]+z[2529]);
assign {c[2531],s[2530]} = (x[2530]+y[2530]+z[2530]);
assign {c[2532],s[2531]} = (x[2531]+y[2531]+z[2531]);
assign {c[2533],s[2532]} = (x[2532]+y[2532]+z[2532]);
assign {c[2534],s[2533]} = (x[2533]+y[2533]+z[2533]);
assign {c[2535],s[2534]} = (x[2534]+y[2534]+z[2534]);
assign {c[2536],s[2535]} = (x[2535]+y[2535]+z[2535]);
assign {c[2537],s[2536]} = (x[2536]+y[2536]+z[2536]);
assign {c[2538],s[2537]} = (x[2537]+y[2537]+z[2537]);
assign {c[2539],s[2538]} = (x[2538]+y[2538]+z[2538]);
assign {c[2540],s[2539]} = (x[2539]+y[2539]+z[2539]);
assign {c[2541],s[2540]} = (x[2540]+y[2540]+z[2540]);
assign {c[2542],s[2541]} = (x[2541]+y[2541]+z[2541]);
assign {c[2543],s[2542]} = (x[2542]+y[2542]+z[2542]);
assign {c[2544],s[2543]} = (x[2543]+y[2543]+z[2543]);
assign {c[2545],s[2544]} = (x[2544]+y[2544]+z[2544]);
assign {c[2546],s[2545]} = (x[2545]+y[2545]+z[2545]);
assign {c[2547],s[2546]} = (x[2546]+y[2546]+z[2546]);
assign {c[2548],s[2547]} = (x[2547]+y[2547]+z[2547]);
assign {c[2549],s[2548]} = (x[2548]+y[2548]+z[2548]);
assign {c[2550],s[2549]} = (x[2549]+y[2549]+z[2549]);
assign {c[2551],s[2550]} = (x[2550]+y[2550]+z[2550]);
assign {c[2552],s[2551]} = (x[2551]+y[2551]+z[2551]);
assign {c[2553],s[2552]} = (x[2552]+y[2552]+z[2552]);
assign {c[2554],s[2553]} = (x[2553]+y[2553]+z[2553]);
assign {c[2555],s[2554]} = (x[2554]+y[2554]+z[2554]);
assign {c[2556],s[2555]} = (x[2555]+y[2555]+z[2555]);
assign {c[2557],s[2556]} = (x[2556]+y[2556]+z[2556]);
assign {c[2558],s[2557]} = (x[2557]+y[2557]+z[2557]);
assign {c[2559],s[2558]} = (x[2558]+y[2558]+z[2558]);
assign {c[2560],s[2559]} = (x[2559]+y[2559]+z[2559]);
assign {c[2561],s[2560]} = (x[2560]+y[2560]+z[2560]);
assign {c[2562],s[2561]} = (x[2561]+y[2561]+z[2561]);
assign {c[2563],s[2562]} = (x[2562]+y[2562]+z[2562]);
assign {c[2564],s[2563]} = (x[2563]+y[2563]+z[2563]);
assign {c[2565],s[2564]} = (x[2564]+y[2564]+z[2564]);
assign {c[2566],s[2565]} = (x[2565]+y[2565]+z[2565]);
assign {c[2567],s[2566]} = (x[2566]+y[2566]+z[2566]);
assign {c[2568],s[2567]} = (x[2567]+y[2567]+z[2567]);
assign {c[2569],s[2568]} = (x[2568]+y[2568]+z[2568]);
assign {c[2570],s[2569]} = (x[2569]+y[2569]+z[2569]);
assign {c[2571],s[2570]} = (x[2570]+y[2570]+z[2570]);
assign {c[2572],s[2571]} = (x[2571]+y[2571]+z[2571]);
assign {c[2573],s[2572]} = (x[2572]+y[2572]+z[2572]);
assign {c[2574],s[2573]} = (x[2573]+y[2573]+z[2573]);
assign {c[2575],s[2574]} = (x[2574]+y[2574]+z[2574]);
assign {c[2576],s[2575]} = (x[2575]+y[2575]+z[2575]);
assign {c[2577],s[2576]} = (x[2576]+y[2576]+z[2576]);
assign {c[2578],s[2577]} = (x[2577]+y[2577]+z[2577]);
assign {c[2579],s[2578]} = (x[2578]+y[2578]+z[2578]);
assign {c[2580],s[2579]} = (x[2579]+y[2579]+z[2579]);
assign {c[2581],s[2580]} = (x[2580]+y[2580]+z[2580]);
assign {c[2582],s[2581]} = (x[2581]+y[2581]+z[2581]);
assign {c[2583],s[2582]} = (x[2582]+y[2582]+z[2582]);
assign {c[2584],s[2583]} = (x[2583]+y[2583]+z[2583]);
assign {c[2585],s[2584]} = (x[2584]+y[2584]+z[2584]);
assign {c[2586],s[2585]} = (x[2585]+y[2585]+z[2585]);
assign {c[2587],s[2586]} = (x[2586]+y[2586]+z[2586]);
assign {c[2588],s[2587]} = (x[2587]+y[2587]+z[2587]);
assign {c[2589],s[2588]} = (x[2588]+y[2588]+z[2588]);
assign {c[2590],s[2589]} = (x[2589]+y[2589]+z[2589]);
assign {c[2591],s[2590]} = (x[2590]+y[2590]+z[2590]);
assign {c[2592],s[2591]} = (x[2591]+y[2591]+z[2591]);
assign {c[2593],s[2592]} = (x[2592]+y[2592]+z[2592]);
assign {c[2594],s[2593]} = (x[2593]+y[2593]+z[2593]);
assign {c[2595],s[2594]} = (x[2594]+y[2594]+z[2594]);
assign {c[2596],s[2595]} = (x[2595]+y[2595]+z[2595]);
assign {c[2597],s[2596]} = (x[2596]+y[2596]+z[2596]);
assign {c[2598],s[2597]} = (x[2597]+y[2597]+z[2597]);
assign {c[2599],s[2598]} = (x[2598]+y[2598]+z[2598]);
assign {c[2600],s[2599]} = (x[2599]+y[2599]+z[2599]);
assign {c[2601],s[2600]} = (x[2600]+y[2600]+z[2600]);
assign {c[2602],s[2601]} = (x[2601]+y[2601]+z[2601]);
assign {c[2603],s[2602]} = (x[2602]+y[2602]+z[2602]);
assign {c[2604],s[2603]} = (x[2603]+y[2603]+z[2603]);
assign {c[2605],s[2604]} = (x[2604]+y[2604]+z[2604]);
assign {c[2606],s[2605]} = (x[2605]+y[2605]+z[2605]);
assign {c[2607],s[2606]} = (x[2606]+y[2606]+z[2606]);
assign {c[2608],s[2607]} = (x[2607]+y[2607]+z[2607]);
assign {c[2609],s[2608]} = (x[2608]+y[2608]+z[2608]);
assign {c[2610],s[2609]} = (x[2609]+y[2609]+z[2609]);
assign {c[2611],s[2610]} = (x[2610]+y[2610]+z[2610]);
assign {c[2612],s[2611]} = (x[2611]+y[2611]+z[2611]);
assign {c[2613],s[2612]} = (x[2612]+y[2612]+z[2612]);
assign {c[2614],s[2613]} = (x[2613]+y[2613]+z[2613]);
assign {c[2615],s[2614]} = (x[2614]+y[2614]+z[2614]);
assign {c[2616],s[2615]} = (x[2615]+y[2615]+z[2615]);
assign {c[2617],s[2616]} = (x[2616]+y[2616]+z[2616]);
assign {c[2618],s[2617]} = (x[2617]+y[2617]+z[2617]);
assign {c[2619],s[2618]} = (x[2618]+y[2618]+z[2618]);
assign {c[2620],s[2619]} = (x[2619]+y[2619]+z[2619]);
assign {c[2621],s[2620]} = (x[2620]+y[2620]+z[2620]);
assign {c[2622],s[2621]} = (x[2621]+y[2621]+z[2621]);
assign {c[2623],s[2622]} = (x[2622]+y[2622]+z[2622]);
assign {c[2624],s[2623]} = (x[2623]+y[2623]+z[2623]);
assign {c[2625],s[2624]} = (x[2624]+y[2624]+z[2624]);
assign {c[2626],s[2625]} = (x[2625]+y[2625]+z[2625]);
assign {c[2627],s[2626]} = (x[2626]+y[2626]+z[2626]);
assign {c[2628],s[2627]} = (x[2627]+y[2627]+z[2627]);
assign {c[2629],s[2628]} = (x[2628]+y[2628]+z[2628]);
assign {c[2630],s[2629]} = (x[2629]+y[2629]+z[2629]);
assign {c[2631],s[2630]} = (x[2630]+y[2630]+z[2630]);
assign {c[2632],s[2631]} = (x[2631]+y[2631]+z[2631]);
assign {c[2633],s[2632]} = (x[2632]+y[2632]+z[2632]);
assign {c[2634],s[2633]} = (x[2633]+y[2633]+z[2633]);
assign {c[2635],s[2634]} = (x[2634]+y[2634]+z[2634]);
assign {c[2636],s[2635]} = (x[2635]+y[2635]+z[2635]);
assign {c[2637],s[2636]} = (x[2636]+y[2636]+z[2636]);
assign {c[2638],s[2637]} = (x[2637]+y[2637]+z[2637]);
assign {c[2639],s[2638]} = (x[2638]+y[2638]+z[2638]);
assign {c[2640],s[2639]} = (x[2639]+y[2639]+z[2639]);
assign {c[2641],s[2640]} = (x[2640]+y[2640]+z[2640]);
assign {c[2642],s[2641]} = (x[2641]+y[2641]+z[2641]);
assign {c[2643],s[2642]} = (x[2642]+y[2642]+z[2642]);
assign {c[2644],s[2643]} = (x[2643]+y[2643]+z[2643]);
assign {c[2645],s[2644]} = (x[2644]+y[2644]+z[2644]);
assign {c[2646],s[2645]} = (x[2645]+y[2645]+z[2645]);
assign {c[2647],s[2646]} = (x[2646]+y[2646]+z[2646]);
assign {c[2648],s[2647]} = (x[2647]+y[2647]+z[2647]);
assign {c[2649],s[2648]} = (x[2648]+y[2648]+z[2648]);
assign {c[2650],s[2649]} = (x[2649]+y[2649]+z[2649]);
assign {c[2651],s[2650]} = (x[2650]+y[2650]+z[2650]);
assign {c[2652],s[2651]} = (x[2651]+y[2651]+z[2651]);
assign {c[2653],s[2652]} = (x[2652]+y[2652]+z[2652]);
assign {c[2654],s[2653]} = (x[2653]+y[2653]+z[2653]);
assign {c[2655],s[2654]} = (x[2654]+y[2654]+z[2654]);
assign {c[2656],s[2655]} = (x[2655]+y[2655]+z[2655]);
assign {c[2657],s[2656]} = (x[2656]+y[2656]+z[2656]);
assign {c[2658],s[2657]} = (x[2657]+y[2657]+z[2657]);
assign {c[2659],s[2658]} = (x[2658]+y[2658]+z[2658]);
assign {c[2660],s[2659]} = (x[2659]+y[2659]+z[2659]);
assign {c[2661],s[2660]} = (x[2660]+y[2660]+z[2660]);
assign {c[2662],s[2661]} = (x[2661]+y[2661]+z[2661]);
assign {c[2663],s[2662]} = (x[2662]+y[2662]+z[2662]);
assign {c[2664],s[2663]} = (x[2663]+y[2663]+z[2663]);
assign {c[2665],s[2664]} = (x[2664]+y[2664]+z[2664]);
assign {c[2666],s[2665]} = (x[2665]+y[2665]+z[2665]);
assign {c[2667],s[2666]} = (x[2666]+y[2666]+z[2666]);
assign {c[2668],s[2667]} = (x[2667]+y[2667]+z[2667]);
assign {c[2669],s[2668]} = (x[2668]+y[2668]+z[2668]);
assign {c[2670],s[2669]} = (x[2669]+y[2669]+z[2669]);
assign {c[2671],s[2670]} = (x[2670]+y[2670]+z[2670]);
assign {c[2672],s[2671]} = (x[2671]+y[2671]+z[2671]);
assign {c[2673],s[2672]} = (x[2672]+y[2672]+z[2672]);
assign {c[2674],s[2673]} = (x[2673]+y[2673]+z[2673]);
assign {c[2675],s[2674]} = (x[2674]+y[2674]+z[2674]);
assign {c[2676],s[2675]} = (x[2675]+y[2675]+z[2675]);
assign {c[2677],s[2676]} = (x[2676]+y[2676]+z[2676]);
assign {c[2678],s[2677]} = (x[2677]+y[2677]+z[2677]);
assign {c[2679],s[2678]} = (x[2678]+y[2678]+z[2678]);
assign {c[2680],s[2679]} = (x[2679]+y[2679]+z[2679]);
assign {c[2681],s[2680]} = (x[2680]+y[2680]+z[2680]);
assign {c[2682],s[2681]} = (x[2681]+y[2681]+z[2681]);
assign {c[2683],s[2682]} = (x[2682]+y[2682]+z[2682]);
assign {c[2684],s[2683]} = (x[2683]+y[2683]+z[2683]);
assign {c[2685],s[2684]} = (x[2684]+y[2684]+z[2684]);
assign {c[2686],s[2685]} = (x[2685]+y[2685]+z[2685]);
assign {c[2687],s[2686]} = (x[2686]+y[2686]+z[2686]);
assign {c[2688],s[2687]} = (x[2687]+y[2687]+z[2687]);
assign {c[2689],s[2688]} = (x[2688]+y[2688]+z[2688]);
assign {c[2690],s[2689]} = (x[2689]+y[2689]+z[2689]);
assign {c[2691],s[2690]} = (x[2690]+y[2690]+z[2690]);
assign {c[2692],s[2691]} = (x[2691]+y[2691]+z[2691]);
assign {c[2693],s[2692]} = (x[2692]+y[2692]+z[2692]);
assign {c[2694],s[2693]} = (x[2693]+y[2693]+z[2693]);
assign {c[2695],s[2694]} = (x[2694]+y[2694]+z[2694]);
assign {c[2696],s[2695]} = (x[2695]+y[2695]+z[2695]);
assign {c[2697],s[2696]} = (x[2696]+y[2696]+z[2696]);
assign {c[2698],s[2697]} = (x[2697]+y[2697]+z[2697]);
assign {c[2699],s[2698]} = (x[2698]+y[2698]+z[2698]);
assign {c[2700],s[2699]} = (x[2699]+y[2699]+z[2699]);
assign {c[2701],s[2700]} = (x[2700]+y[2700]+z[2700]);
assign {c[2702],s[2701]} = (x[2701]+y[2701]+z[2701]);
assign {c[2703],s[2702]} = (x[2702]+y[2702]+z[2702]);
assign {c[2704],s[2703]} = (x[2703]+y[2703]+z[2703]);
assign {c[2705],s[2704]} = (x[2704]+y[2704]+z[2704]);
assign {c[2706],s[2705]} = (x[2705]+y[2705]+z[2705]);
assign {c[2707],s[2706]} = (x[2706]+y[2706]+z[2706]);
assign {c[2708],s[2707]} = (x[2707]+y[2707]+z[2707]);
assign {c[2709],s[2708]} = (x[2708]+y[2708]+z[2708]);
assign {c[2710],s[2709]} = (x[2709]+y[2709]+z[2709]);
assign {c[2711],s[2710]} = (x[2710]+y[2710]+z[2710]);
assign {c[2712],s[2711]} = (x[2711]+y[2711]+z[2711]);
assign {c[2713],s[2712]} = (x[2712]+y[2712]+z[2712]);
assign {c[2714],s[2713]} = (x[2713]+y[2713]+z[2713]);
assign {c[2715],s[2714]} = (x[2714]+y[2714]+z[2714]);
assign {c[2716],s[2715]} = (x[2715]+y[2715]+z[2715]);
assign {c[2717],s[2716]} = (x[2716]+y[2716]+z[2716]);
assign {c[2718],s[2717]} = (x[2717]+y[2717]+z[2717]);
assign {c[2719],s[2718]} = (x[2718]+y[2718]+z[2718]);
assign {c[2720],s[2719]} = (x[2719]+y[2719]+z[2719]);
assign {c[2721],s[2720]} = (x[2720]+y[2720]+z[2720]);
assign {c[2722],s[2721]} = (x[2721]+y[2721]+z[2721]);
assign {c[2723],s[2722]} = (x[2722]+y[2722]+z[2722]);
assign {c[2724],s[2723]} = (x[2723]+y[2723]+z[2723]);
assign {c[2725],s[2724]} = (x[2724]+y[2724]+z[2724]);
assign {c[2726],s[2725]} = (x[2725]+y[2725]+z[2725]);
assign {c[2727],s[2726]} = (x[2726]+y[2726]+z[2726]);
assign {c[2728],s[2727]} = (x[2727]+y[2727]+z[2727]);
assign {c[2729],s[2728]} = (x[2728]+y[2728]+z[2728]);
assign {c[2730],s[2729]} = (x[2729]+y[2729]+z[2729]);
assign {c[2731],s[2730]} = (x[2730]+y[2730]+z[2730]);
assign {c[2732],s[2731]} = (x[2731]+y[2731]+z[2731]);
assign {c[2733],s[2732]} = (x[2732]+y[2732]+z[2732]);
assign {c[2734],s[2733]} = (x[2733]+y[2733]+z[2733]);
assign {c[2735],s[2734]} = (x[2734]+y[2734]+z[2734]);
assign {c[2736],s[2735]} = (x[2735]+y[2735]+z[2735]);
assign {c[2737],s[2736]} = (x[2736]+y[2736]+z[2736]);
assign {c[2738],s[2737]} = (x[2737]+y[2737]+z[2737]);
assign {c[2739],s[2738]} = (x[2738]+y[2738]+z[2738]);
assign {c[2740],s[2739]} = (x[2739]+y[2739]+z[2739]);
assign {c[2741],s[2740]} = (x[2740]+y[2740]+z[2740]);
assign {c[2742],s[2741]} = (x[2741]+y[2741]+z[2741]);
assign {c[2743],s[2742]} = (x[2742]+y[2742]+z[2742]);
assign {c[2744],s[2743]} = (x[2743]+y[2743]+z[2743]);
assign {c[2745],s[2744]} = (x[2744]+y[2744]+z[2744]);
assign {c[2746],s[2745]} = (x[2745]+y[2745]+z[2745]);
assign {c[2747],s[2746]} = (x[2746]+y[2746]+z[2746]);
assign {c[2748],s[2747]} = (x[2747]+y[2747]+z[2747]);
assign {c[2749],s[2748]} = (x[2748]+y[2748]+z[2748]);
assign {c[2750],s[2749]} = (x[2749]+y[2749]+z[2749]);
assign {c[2751],s[2750]} = (x[2750]+y[2750]+z[2750]);
assign {c[2752],s[2751]} = (x[2751]+y[2751]+z[2751]);
assign {c[2753],s[2752]} = (x[2752]+y[2752]+z[2752]);
assign {c[2754],s[2753]} = (x[2753]+y[2753]+z[2753]);
assign {c[2755],s[2754]} = (x[2754]+y[2754]+z[2754]);
assign {c[2756],s[2755]} = (x[2755]+y[2755]+z[2755]);
assign {c[2757],s[2756]} = (x[2756]+y[2756]+z[2756]);
assign {c[2758],s[2757]} = (x[2757]+y[2757]+z[2757]);
assign {c[2759],s[2758]} = (x[2758]+y[2758]+z[2758]);
assign {c[2760],s[2759]} = (x[2759]+y[2759]+z[2759]);
assign {c[2761],s[2760]} = (x[2760]+y[2760]+z[2760]);
assign {c[2762],s[2761]} = (x[2761]+y[2761]+z[2761]);
assign {c[2763],s[2762]} = (x[2762]+y[2762]+z[2762]);
assign {c[2764],s[2763]} = (x[2763]+y[2763]+z[2763]);
assign {c[2765],s[2764]} = (x[2764]+y[2764]+z[2764]);
assign {c[2766],s[2765]} = (x[2765]+y[2765]+z[2765]);
assign {c[2767],s[2766]} = (x[2766]+y[2766]+z[2766]);
assign {c[2768],s[2767]} = (x[2767]+y[2767]+z[2767]);
assign {c[2769],s[2768]} = (x[2768]+y[2768]+z[2768]);
assign {c[2770],s[2769]} = (x[2769]+y[2769]+z[2769]);
assign {c[2771],s[2770]} = (x[2770]+y[2770]+z[2770]);
assign {c[2772],s[2771]} = (x[2771]+y[2771]+z[2771]);
assign {c[2773],s[2772]} = (x[2772]+y[2772]+z[2772]);
assign {c[2774],s[2773]} = (x[2773]+y[2773]+z[2773]);
assign {c[2775],s[2774]} = (x[2774]+y[2774]+z[2774]);
assign {c[2776],s[2775]} = (x[2775]+y[2775]+z[2775]);
assign {c[2777],s[2776]} = (x[2776]+y[2776]+z[2776]);
assign {c[2778],s[2777]} = (x[2777]+y[2777]+z[2777]);
assign {c[2779],s[2778]} = (x[2778]+y[2778]+z[2778]);
assign {c[2780],s[2779]} = (x[2779]+y[2779]+z[2779]);
assign {c[2781],s[2780]} = (x[2780]+y[2780]+z[2780]);
assign {c[2782],s[2781]} = (x[2781]+y[2781]+z[2781]);
assign {c[2783],s[2782]} = (x[2782]+y[2782]+z[2782]);
assign {c[2784],s[2783]} = (x[2783]+y[2783]+z[2783]);
assign {c[2785],s[2784]} = (x[2784]+y[2784]+z[2784]);
assign {c[2786],s[2785]} = (x[2785]+y[2785]+z[2785]);
assign {c[2787],s[2786]} = (x[2786]+y[2786]+z[2786]);
assign {c[2788],s[2787]} = (x[2787]+y[2787]+z[2787]);
assign {c[2789],s[2788]} = (x[2788]+y[2788]+z[2788]);
assign {c[2790],s[2789]} = (x[2789]+y[2789]+z[2789]);
assign {c[2791],s[2790]} = (x[2790]+y[2790]+z[2790]);
assign {c[2792],s[2791]} = (x[2791]+y[2791]+z[2791]);
assign {c[2793],s[2792]} = (x[2792]+y[2792]+z[2792]);
assign {c[2794],s[2793]} = (x[2793]+y[2793]+z[2793]);
assign {c[2795],s[2794]} = (x[2794]+y[2794]+z[2794]);
assign {c[2796],s[2795]} = (x[2795]+y[2795]+z[2795]);
assign {c[2797],s[2796]} = (x[2796]+y[2796]+z[2796]);
assign {c[2798],s[2797]} = (x[2797]+y[2797]+z[2797]);
assign {c[2799],s[2798]} = (x[2798]+y[2798]+z[2798]);
assign {c[2800],s[2799]} = (x[2799]+y[2799]+z[2799]);
assign {c[2801],s[2800]} = (x[2800]+y[2800]+z[2800]);
assign {c[2802],s[2801]} = (x[2801]+y[2801]+z[2801]);
assign {c[2803],s[2802]} = (x[2802]+y[2802]+z[2802]);
assign {c[2804],s[2803]} = (x[2803]+y[2803]+z[2803]);
assign {c[2805],s[2804]} = (x[2804]+y[2804]+z[2804]);
assign {c[2806],s[2805]} = (x[2805]+y[2805]+z[2805]);
assign {c[2807],s[2806]} = (x[2806]+y[2806]+z[2806]);
assign {c[2808],s[2807]} = (x[2807]+y[2807]+z[2807]);
assign {c[2809],s[2808]} = (x[2808]+y[2808]+z[2808]);
assign {c[2810],s[2809]} = (x[2809]+y[2809]+z[2809]);
assign {c[2811],s[2810]} = (x[2810]+y[2810]+z[2810]);
assign {c[2812],s[2811]} = (x[2811]+y[2811]+z[2811]);
assign {c[2813],s[2812]} = (x[2812]+y[2812]+z[2812]);
assign {c[2814],s[2813]} = (x[2813]+y[2813]+z[2813]);
assign {c[2815],s[2814]} = (x[2814]+y[2814]+z[2814]);
assign {c[2816],s[2815]} = (x[2815]+y[2815]+z[2815]);
assign {c[2817],s[2816]} = (x[2816]+y[2816]+z[2816]);
assign {c[2818],s[2817]} = (x[2817]+y[2817]+z[2817]);
assign {c[2819],s[2818]} = (x[2818]+y[2818]+z[2818]);
assign {c[2820],s[2819]} = (x[2819]+y[2819]+z[2819]);
assign {c[2821],s[2820]} = (x[2820]+y[2820]+z[2820]);
assign {c[2822],s[2821]} = (x[2821]+y[2821]+z[2821]);
assign {c[2823],s[2822]} = (x[2822]+y[2822]+z[2822]);
assign {c[2824],s[2823]} = (x[2823]+y[2823]+z[2823]);
assign {c[2825],s[2824]} = (x[2824]+y[2824]+z[2824]);
assign {c[2826],s[2825]} = (x[2825]+y[2825]+z[2825]);
assign {c[2827],s[2826]} = (x[2826]+y[2826]+z[2826]);
assign {c[2828],s[2827]} = (x[2827]+y[2827]+z[2827]);
assign {c[2829],s[2828]} = (x[2828]+y[2828]+z[2828]);
assign {c[2830],s[2829]} = (x[2829]+y[2829]+z[2829]);
assign {c[2831],s[2830]} = (x[2830]+y[2830]+z[2830]);
assign {c[2832],s[2831]} = (x[2831]+y[2831]+z[2831]);
assign {c[2833],s[2832]} = (x[2832]+y[2832]+z[2832]);
assign {c[2834],s[2833]} = (x[2833]+y[2833]+z[2833]);
assign {c[2835],s[2834]} = (x[2834]+y[2834]+z[2834]);
assign {c[2836],s[2835]} = (x[2835]+y[2835]+z[2835]);
assign {c[2837],s[2836]} = (x[2836]+y[2836]+z[2836]);
assign {c[2838],s[2837]} = (x[2837]+y[2837]+z[2837]);
assign {c[2839],s[2838]} = (x[2838]+y[2838]+z[2838]);
assign {c[2840],s[2839]} = (x[2839]+y[2839]+z[2839]);
assign {c[2841],s[2840]} = (x[2840]+y[2840]+z[2840]);
assign {c[2842],s[2841]} = (x[2841]+y[2841]+z[2841]);
assign {c[2843],s[2842]} = (x[2842]+y[2842]+z[2842]);
assign {c[2844],s[2843]} = (x[2843]+y[2843]+z[2843]);
assign {c[2845],s[2844]} = (x[2844]+y[2844]+z[2844]);
assign {c[2846],s[2845]} = (x[2845]+y[2845]+z[2845]);
assign {c[2847],s[2846]} = (x[2846]+y[2846]+z[2846]);
assign {c[2848],s[2847]} = (x[2847]+y[2847]+z[2847]);
assign {c[2849],s[2848]} = (x[2848]+y[2848]+z[2848]);
assign {c[2850],s[2849]} = (x[2849]+y[2849]+z[2849]);
assign {c[2851],s[2850]} = (x[2850]+y[2850]+z[2850]);
assign {c[2852],s[2851]} = (x[2851]+y[2851]+z[2851]);
assign {c[2853],s[2852]} = (x[2852]+y[2852]+z[2852]);
assign {c[2854],s[2853]} = (x[2853]+y[2853]+z[2853]);
assign {c[2855],s[2854]} = (x[2854]+y[2854]+z[2854]);
assign {c[2856],s[2855]} = (x[2855]+y[2855]+z[2855]);
assign {c[2857],s[2856]} = (x[2856]+y[2856]+z[2856]);
assign {c[2858],s[2857]} = (x[2857]+y[2857]+z[2857]);
assign {c[2859],s[2858]} = (x[2858]+y[2858]+z[2858]);
assign {c[2860],s[2859]} = (x[2859]+y[2859]+z[2859]);
assign {c[2861],s[2860]} = (x[2860]+y[2860]+z[2860]);
assign {c[2862],s[2861]} = (x[2861]+y[2861]+z[2861]);
assign {c[2863],s[2862]} = (x[2862]+y[2862]+z[2862]);
assign {c[2864],s[2863]} = (x[2863]+y[2863]+z[2863]);
assign {c[2865],s[2864]} = (x[2864]+y[2864]+z[2864]);
assign {c[2866],s[2865]} = (x[2865]+y[2865]+z[2865]);
assign {c[2867],s[2866]} = (x[2866]+y[2866]+z[2866]);
assign {c[2868],s[2867]} = (x[2867]+y[2867]+z[2867]);
assign {c[2869],s[2868]} = (x[2868]+y[2868]+z[2868]);
assign {c[2870],s[2869]} = (x[2869]+y[2869]+z[2869]);
assign {c[2871],s[2870]} = (x[2870]+y[2870]+z[2870]);
assign {c[2872],s[2871]} = (x[2871]+y[2871]+z[2871]);
assign {c[2873],s[2872]} = (x[2872]+y[2872]+z[2872]);
assign {c[2874],s[2873]} = (x[2873]+y[2873]+z[2873]);
assign {c[2875],s[2874]} = (x[2874]+y[2874]+z[2874]);
assign {c[2876],s[2875]} = (x[2875]+y[2875]+z[2875]);
assign {c[2877],s[2876]} = (x[2876]+y[2876]+z[2876]);
assign {c[2878],s[2877]} = (x[2877]+y[2877]+z[2877]);
assign {c[2879],s[2878]} = (x[2878]+y[2878]+z[2878]);
assign {c[2880],s[2879]} = (x[2879]+y[2879]+z[2879]);
assign {c[2881],s[2880]} = (x[2880]+y[2880]+z[2880]);
assign {c[2882],s[2881]} = (x[2881]+y[2881]+z[2881]);
assign {c[2883],s[2882]} = (x[2882]+y[2882]+z[2882]);
assign {c[2884],s[2883]} = (x[2883]+y[2883]+z[2883]);
assign {c[2885],s[2884]} = (x[2884]+y[2884]+z[2884]);
assign {c[2886],s[2885]} = (x[2885]+y[2885]+z[2885]);
assign {c[2887],s[2886]} = (x[2886]+y[2886]+z[2886]);
assign {c[2888],s[2887]} = (x[2887]+y[2887]+z[2887]);
assign {c[2889],s[2888]} = (x[2888]+y[2888]+z[2888]);
assign {c[2890],s[2889]} = (x[2889]+y[2889]+z[2889]);
assign {c[2891],s[2890]} = (x[2890]+y[2890]+z[2890]);
assign {c[2892],s[2891]} = (x[2891]+y[2891]+z[2891]);
assign {c[2893],s[2892]} = (x[2892]+y[2892]+z[2892]);
assign {c[2894],s[2893]} = (x[2893]+y[2893]+z[2893]);
assign {c[2895],s[2894]} = (x[2894]+y[2894]+z[2894]);
assign {c[2896],s[2895]} = (x[2895]+y[2895]+z[2895]);
assign {c[2897],s[2896]} = (x[2896]+y[2896]+z[2896]);
assign {c[2898],s[2897]} = (x[2897]+y[2897]+z[2897]);
assign {c[2899],s[2898]} = (x[2898]+y[2898]+z[2898]);
assign {c[2900],s[2899]} = (x[2899]+y[2899]+z[2899]);
assign {c[2901],s[2900]} = (x[2900]+y[2900]+z[2900]);
assign {c[2902],s[2901]} = (x[2901]+y[2901]+z[2901]);
assign {c[2903],s[2902]} = (x[2902]+y[2902]+z[2902]);
assign {c[2904],s[2903]} = (x[2903]+y[2903]+z[2903]);
assign {c[2905],s[2904]} = (x[2904]+y[2904]+z[2904]);
assign {c[2906],s[2905]} = (x[2905]+y[2905]+z[2905]);
assign {c[2907],s[2906]} = (x[2906]+y[2906]+z[2906]);
assign {c[2908],s[2907]} = (x[2907]+y[2907]+z[2907]);
assign {c[2909],s[2908]} = (x[2908]+y[2908]+z[2908]);
assign {c[2910],s[2909]} = (x[2909]+y[2909]+z[2909]);
assign {c[2911],s[2910]} = (x[2910]+y[2910]+z[2910]);
assign {c[2912],s[2911]} = (x[2911]+y[2911]+z[2911]);
assign {c[2913],s[2912]} = (x[2912]+y[2912]+z[2912]);
assign {c[2914],s[2913]} = (x[2913]+y[2913]+z[2913]);
assign {c[2915],s[2914]} = (x[2914]+y[2914]+z[2914]);
assign {c[2916],s[2915]} = (x[2915]+y[2915]+z[2915]);
assign {c[2917],s[2916]} = (x[2916]+y[2916]+z[2916]);
assign {c[2918],s[2917]} = (x[2917]+y[2917]+z[2917]);
assign {c[2919],s[2918]} = (x[2918]+y[2918]+z[2918]);
assign {c[2920],s[2919]} = (x[2919]+y[2919]+z[2919]);
assign {c[2921],s[2920]} = (x[2920]+y[2920]+z[2920]);
assign {c[2922],s[2921]} = (x[2921]+y[2921]+z[2921]);
assign {c[2923],s[2922]} = (x[2922]+y[2922]+z[2922]);
assign {c[2924],s[2923]} = (x[2923]+y[2923]+z[2923]);
assign {c[2925],s[2924]} = (x[2924]+y[2924]+z[2924]);
assign {c[2926],s[2925]} = (x[2925]+y[2925]+z[2925]);
assign {c[2927],s[2926]} = (x[2926]+y[2926]+z[2926]);
assign {c[2928],s[2927]} = (x[2927]+y[2927]+z[2927]);
assign {c[2929],s[2928]} = (x[2928]+y[2928]+z[2928]);
assign {c[2930],s[2929]} = (x[2929]+y[2929]+z[2929]);
assign {c[2931],s[2930]} = (x[2930]+y[2930]+z[2930]);
assign {c[2932],s[2931]} = (x[2931]+y[2931]+z[2931]);
assign {c[2933],s[2932]} = (x[2932]+y[2932]+z[2932]);
assign {c[2934],s[2933]} = (x[2933]+y[2933]+z[2933]);
assign {c[2935],s[2934]} = (x[2934]+y[2934]+z[2934]);
assign {c[2936],s[2935]} = (x[2935]+y[2935]+z[2935]);
assign {c[2937],s[2936]} = (x[2936]+y[2936]+z[2936]);
assign {c[2938],s[2937]} = (x[2937]+y[2937]+z[2937]);
assign {c[2939],s[2938]} = (x[2938]+y[2938]+z[2938]);
assign {c[2940],s[2939]} = (x[2939]+y[2939]+z[2939]);
assign {c[2941],s[2940]} = (x[2940]+y[2940]+z[2940]);
assign {c[2942],s[2941]} = (x[2941]+y[2941]+z[2941]);
assign {c[2943],s[2942]} = (x[2942]+y[2942]+z[2942]);
assign {c[2944],s[2943]} = (x[2943]+y[2943]+z[2943]);
assign {c[2945],s[2944]} = (x[2944]+y[2944]+z[2944]);
assign {c[2946],s[2945]} = (x[2945]+y[2945]+z[2945]);
assign {c[2947],s[2946]} = (x[2946]+y[2946]+z[2946]);
assign {c[2948],s[2947]} = (x[2947]+y[2947]+z[2947]);
assign {c[2949],s[2948]} = (x[2948]+y[2948]+z[2948]);
assign {c[2950],s[2949]} = (x[2949]+y[2949]+z[2949]);
assign {c[2951],s[2950]} = (x[2950]+y[2950]+z[2950]);
assign {c[2952],s[2951]} = (x[2951]+y[2951]+z[2951]);
assign {c[2953],s[2952]} = (x[2952]+y[2952]+z[2952]);
assign {c[2954],s[2953]} = (x[2953]+y[2953]+z[2953]);
assign {c[2955],s[2954]} = (x[2954]+y[2954]+z[2954]);
assign {c[2956],s[2955]} = (x[2955]+y[2955]+z[2955]);
assign {c[2957],s[2956]} = (x[2956]+y[2956]+z[2956]);
assign {c[2958],s[2957]} = (x[2957]+y[2957]+z[2957]);
assign {c[2959],s[2958]} = (x[2958]+y[2958]+z[2958]);
assign {c[2960],s[2959]} = (x[2959]+y[2959]+z[2959]);
assign {c[2961],s[2960]} = (x[2960]+y[2960]+z[2960]);
assign {c[2962],s[2961]} = (x[2961]+y[2961]+z[2961]);
assign {c[2963],s[2962]} = (x[2962]+y[2962]+z[2962]);
assign {c[2964],s[2963]} = (x[2963]+y[2963]+z[2963]);
assign {c[2965],s[2964]} = (x[2964]+y[2964]+z[2964]);
assign {c[2966],s[2965]} = (x[2965]+y[2965]+z[2965]);
assign {c[2967],s[2966]} = (x[2966]+y[2966]+z[2966]);
assign {c[2968],s[2967]} = (x[2967]+y[2967]+z[2967]);
assign {c[2969],s[2968]} = (x[2968]+y[2968]+z[2968]);
assign {c[2970],s[2969]} = (x[2969]+y[2969]+z[2969]);
assign {c[2971],s[2970]} = (x[2970]+y[2970]+z[2970]);
assign {c[2972],s[2971]} = (x[2971]+y[2971]+z[2971]);
assign {c[2973],s[2972]} = (x[2972]+y[2972]+z[2972]);
assign {c[2974],s[2973]} = (x[2973]+y[2973]+z[2973]);
assign {c[2975],s[2974]} = (x[2974]+y[2974]+z[2974]);
assign {c[2976],s[2975]} = (x[2975]+y[2975]+z[2975]);
assign {c[2977],s[2976]} = (x[2976]+y[2976]+z[2976]);
assign {c[2978],s[2977]} = (x[2977]+y[2977]+z[2977]);
assign {c[2979],s[2978]} = (x[2978]+y[2978]+z[2978]);
assign {c[2980],s[2979]} = (x[2979]+y[2979]+z[2979]);
assign {c[2981],s[2980]} = (x[2980]+y[2980]+z[2980]);
assign {c[2982],s[2981]} = (x[2981]+y[2981]+z[2981]);
assign {c[2983],s[2982]} = (x[2982]+y[2982]+z[2982]);
assign {c[2984],s[2983]} = (x[2983]+y[2983]+z[2983]);
assign {c[2985],s[2984]} = (x[2984]+y[2984]+z[2984]);
assign {c[2986],s[2985]} = (x[2985]+y[2985]+z[2985]);
assign {c[2987],s[2986]} = (x[2986]+y[2986]+z[2986]);
assign {c[2988],s[2987]} = (x[2987]+y[2987]+z[2987]);
assign {c[2989],s[2988]} = (x[2988]+y[2988]+z[2988]);
assign {c[2990],s[2989]} = (x[2989]+y[2989]+z[2989]);
assign {c[2991],s[2990]} = (x[2990]+y[2990]+z[2990]);
assign {c[2992],s[2991]} = (x[2991]+y[2991]+z[2991]);
assign {c[2993],s[2992]} = (x[2992]+y[2992]+z[2992]);
assign {c[2994],s[2993]} = (x[2993]+y[2993]+z[2993]);
assign {c[2995],s[2994]} = (x[2994]+y[2994]+z[2994]);
assign {c[2996],s[2995]} = (x[2995]+y[2995]+z[2995]);
assign {c[2997],s[2996]} = (x[2996]+y[2996]+z[2996]);
assign {c[2998],s[2997]} = (x[2997]+y[2997]+z[2997]);
assign {c[2999],s[2998]} = (x[2998]+y[2998]+z[2998]);
assign {c[3000],s[2999]} = (x[2999]+y[2999]+z[2999]);
assign {c[3001],s[3000]} = (x[3000]+y[3000]+z[3000]);
assign {c[3002],s[3001]} = (x[3001]+y[3001]+z[3001]);
assign {c[3003],s[3002]} = (x[3002]+y[3002]+z[3002]);
assign {c[3004],s[3003]} = (x[3003]+y[3003]+z[3003]);
assign {c[3005],s[3004]} = (x[3004]+y[3004]+z[3004]);
assign {c[3006],s[3005]} = (x[3005]+y[3005]+z[3005]);
assign {c[3007],s[3006]} = (x[3006]+y[3006]+z[3006]);
assign {c[3008],s[3007]} = (x[3007]+y[3007]+z[3007]);
assign {c[3009],s[3008]} = (x[3008]+y[3008]+z[3008]);
assign {c[3010],s[3009]} = (x[3009]+y[3009]+z[3009]);
assign {c[3011],s[3010]} = (x[3010]+y[3010]+z[3010]);
assign {c[3012],s[3011]} = (x[3011]+y[3011]+z[3011]);
assign {c[3013],s[3012]} = (x[3012]+y[3012]+z[3012]);
assign {c[3014],s[3013]} = (x[3013]+y[3013]+z[3013]);
assign {c[3015],s[3014]} = (x[3014]+y[3014]+z[3014]);
assign {c[3016],s[3015]} = (x[3015]+y[3015]+z[3015]);
assign {c[3017],s[3016]} = (x[3016]+y[3016]+z[3016]);
assign {dummy,s[3017]} = (x[3017]+y[3017]+z[3017]);

endmodule
    