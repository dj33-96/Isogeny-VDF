
module AND_matrix_43x43(
    input [42:0] a,
    input [42:0] b,
    output [3697:0] c // lines are appended together
);
    
wire [42:0] c_w_0;
wire [42:0] c_w_1;
wire [42:0] c_w_2;
wire [42:0] c_w_3;
wire [42:0] c_w_4;
wire [42:0] c_w_5;
wire [42:0] c_w_6;
wire [42:0] c_w_7;
wire [42:0] c_w_8;
wire [42:0] c_w_9;
wire [42:0] c_w_10;
wire [42:0] c_w_11;
wire [42:0] c_w_12;
wire [42:0] c_w_13;
wire [42:0] c_w_14;
wire [42:0] c_w_15;
wire [42:0] c_w_16;
wire [42:0] c_w_17;
wire [42:0] c_w_18;
wire [42:0] c_w_19;
wire [42:0] c_w_20;
wire [42:0] c_w_21;
wire [42:0] c_w_22;
wire [42:0] c_w_23;
wire [42:0] c_w_24;
wire [42:0] c_w_25;
wire [42:0] c_w_26;
wire [42:0] c_w_27;
wire [42:0] c_w_28;
wire [42:0] c_w_29;
wire [42:0] c_w_30;
wire [42:0] c_w_31;
wire [42:0] c_w_32;
wire [42:0] c_w_33;
wire [42:0] c_w_34;
wire [42:0] c_w_35;
wire [42:0] c_w_36;
wire [42:0] c_w_37;
wire [42:0] c_w_38;
wire [42:0] c_w_39;
wire [42:0] c_w_40;
wire [42:0] c_w_41;
wire [42:0] c_w_42;
    
AND_array_43 AND_array_43_i0(a,b[0],c_w_0);
AND_array_43 AND_array_43_i1(a,b[1],c_w_1);
AND_array_43 AND_array_43_i2(a,b[2],c_w_2);
AND_array_43 AND_array_43_i3(a,b[3],c_w_3);
AND_array_43 AND_array_43_i4(a,b[4],c_w_4);
AND_array_43 AND_array_43_i5(a,b[5],c_w_5);
AND_array_43 AND_array_43_i6(a,b[6],c_w_6);
AND_array_43 AND_array_43_i7(a,b[7],c_w_7);
AND_array_43 AND_array_43_i8(a,b[8],c_w_8);
AND_array_43 AND_array_43_i9(a,b[9],c_w_9);
AND_array_43 AND_array_43_i10(a,b[10],c_w_10);
AND_array_43 AND_array_43_i11(a,b[11],c_w_11);
AND_array_43 AND_array_43_i12(a,b[12],c_w_12);
AND_array_43 AND_array_43_i13(a,b[13],c_w_13);
AND_array_43 AND_array_43_i14(a,b[14],c_w_14);
AND_array_43 AND_array_43_i15(a,b[15],c_w_15);
AND_array_43 AND_array_43_i16(a,b[16],c_w_16);
AND_array_43 AND_array_43_i17(a,b[17],c_w_17);
AND_array_43 AND_array_43_i18(a,b[18],c_w_18);
AND_array_43 AND_array_43_i19(a,b[19],c_w_19);
AND_array_43 AND_array_43_i20(a,b[20],c_w_20);
AND_array_43 AND_array_43_i21(a,b[21],c_w_21);
AND_array_43 AND_array_43_i22(a,b[22],c_w_22);
AND_array_43 AND_array_43_i23(a,b[23],c_w_23);
AND_array_43 AND_array_43_i24(a,b[24],c_w_24);
AND_array_43 AND_array_43_i25(a,b[25],c_w_25);
AND_array_43 AND_array_43_i26(a,b[26],c_w_26);
AND_array_43 AND_array_43_i27(a,b[27],c_w_27);
AND_array_43 AND_array_43_i28(a,b[28],c_w_28);
AND_array_43 AND_array_43_i29(a,b[29],c_w_29);
AND_array_43 AND_array_43_i30(a,b[30],c_w_30);
AND_array_43 AND_array_43_i31(a,b[31],c_w_31);
AND_array_43 AND_array_43_i32(a,b[32],c_w_32);
AND_array_43 AND_array_43_i33(a,b[33],c_w_33);
AND_array_43 AND_array_43_i34(a,b[34],c_w_34);
AND_array_43 AND_array_43_i35(a,b[35],c_w_35);
AND_array_43 AND_array_43_i36(a,b[36],c_w_36);
AND_array_43 AND_array_43_i37(a,b[37],c_w_37);
AND_array_43 AND_array_43_i38(a,b[38],c_w_38);
AND_array_43 AND_array_43_i39(a,b[39],c_w_39);
AND_array_43 AND_array_43_i40(a,b[40],c_w_40);
AND_array_43 AND_array_43_i41(a,b[41],c_w_41);
AND_array_43 AND_array_43_i42(a,b[42],c_w_42);
    
assign c[85:0] = {43'b0,c_w_0};
assign c[171:86] = {42'b0,c_w_1,1'b0};
assign c[257:172] = {41'b0,c_w_2,2'b0};
assign c[343:258] = {40'b0,c_w_3,3'b0};
assign c[429:344] = {39'b0,c_w_4,4'b0};
assign c[515:430] = {38'b0,c_w_5,5'b0};
assign c[601:516] = {37'b0,c_w_6,6'b0};
assign c[687:602] = {36'b0,c_w_7,7'b0};
assign c[773:688] = {35'b0,c_w_8,8'b0};
assign c[859:774] = {34'b0,c_w_9,9'b0};
assign c[945:860] = {33'b0,c_w_10,10'b0};
assign c[1031:946] = {32'b0,c_w_11,11'b0};
assign c[1117:1032] = {31'b0,c_w_12,12'b0};
assign c[1203:1118] = {30'b0,c_w_13,13'b0};
assign c[1289:1204] = {29'b0,c_w_14,14'b0};
assign c[1375:1290] = {28'b0,c_w_15,15'b0};
assign c[1461:1376] = {27'b0,c_w_16,16'b0};
assign c[1547:1462] = {26'b0,c_w_17,17'b0};
assign c[1633:1548] = {25'b0,c_w_18,18'b0};
assign c[1719:1634] = {24'b0,c_w_19,19'b0};
assign c[1805:1720] = {23'b0,c_w_20,20'b0};
assign c[1891:1806] = {22'b0,c_w_21,21'b0};
assign c[1977:1892] = {21'b0,c_w_22,22'b0};
assign c[2063:1978] = {20'b0,c_w_23,23'b0};
assign c[2149:2064] = {19'b0,c_w_24,24'b0};
assign c[2235:2150] = {18'b0,c_w_25,25'b0};
assign c[2321:2236] = {17'b0,c_w_26,26'b0};
assign c[2407:2322] = {16'b0,c_w_27,27'b0};
assign c[2493:2408] = {15'b0,c_w_28,28'b0};
assign c[2579:2494] = {14'b0,c_w_29,29'b0};
assign c[2665:2580] = {13'b0,c_w_30,30'b0};
assign c[2751:2666] = {12'b0,c_w_31,31'b0};
assign c[2837:2752] = {11'b0,c_w_32,32'b0};
assign c[2923:2838] = {10'b0,c_w_33,33'b0};
assign c[3009:2924] = {9'b0,c_w_34,34'b0};
assign c[3095:3010] = {8'b0,c_w_35,35'b0};
assign c[3181:3096] = {7'b0,c_w_36,36'b0};
assign c[3267:3182] = {6'b0,c_w_37,37'b0};
assign c[3353:3268] = {5'b0,c_w_38,38'b0};
assign c[3439:3354] = {4'b0,c_w_39,39'b0};
assign c[3525:3440] = {3'b0,c_w_40,40'b0};
assign c[3611:3526] = {2'b0,c_w_41,41'b0};
assign c[3697:3612] = {1'b0,c_w_42,42'b0};
    
endmodule
    