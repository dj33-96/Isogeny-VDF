
module ha(
    input x,y,
    output c,s
);

assign {c,s} = x+y;

endmodule
    