
module tb_4_iso_e_1506();

// Instruction list + effect:
/*
INS = 0 => Idle
INS = 1 => load input
INS = 2 => copy point rd to wr
INS = 3 => ADD
INS = 4 => SUB
INS = 5 => MUL
*/

reg clk,rst,get_output,data_en,ins_in;
wire [24-1:0] command_in;
reg [1506-1:0] din_1,din_2;
wire [1506-1:0] dout_1,dout_2;

reg [2:0] INS;
reg [7-1:0] rd_addr_1,rd_addr_2,wr_addr;

assign command_in = {INS,rd_addr_1,rd_addr_2,wr_addr};

wire [1506:0] p, calculated;
assign p = 1507'd1658539334852043956605014686969369842243820155059458240864380460354175875596746126442552006529285980003318752448184629099761975446397870870332614114924526019655624366944770281974501212314250998405682106067115619475132937730960746637418716661215852316737808364060021400361715167852784987427099666051667608448888314571788638487985846716927693574019769274326804364407638203115258648742883949562283207610572974523311143132532016594886767069744238342663307263;
assign calculated = (dout_1 + dout_2) % p;

wire [1506-1:0] x,z,k1,k2,k3;//inputs
wire [1506-1:0] xo,zo;//expected values

assign x = 1506'd1533910757811517331179909129660025853084150426833233172483140215941333894701571607724163540785617560561908071475391513249074982833758318480567484410558066725638717760519355558111099758161765145631561659544230868661091402658244484215666523994536888718591040720663254029460682567379006992919158917480697629007998756326495938081292384853430180689238866059705385770531065903961227622528967924509814888658798393796944939677441028446770220654996788482357298557;
assign z = 1506'd778780221328586877322847292786807663188759349688439660564284398558774481443019423422328877131584858315445859782594757424171559081012287741646926741246683190316977667329522920783653622450509040453386279276466177597905935915139613341954858094088208364530489330988946866583939187786457633569793857674778799530264883305287560334606324370848446108940086367361522458058491233628818600600584037346745976236507207103989127465641762293773048958642348525650191515;
assign k1 = 1506'd632488848111606046430876648175092098662326213823486762189754012090936105036496993596844713019145766044046054941703471611534442768354210373002201448332957499112142275497209922238593633285536842001877321699824749819728280810961038537070541159555638775796098575567291548980439938438659294495864071689849582809414400570077775229255036986797066525436158054446621297898177119819100299379235975937584080315844958490488476474218765956830785876051293242157221353;
assign k2 = 1506'd696318202978316488695558868226104574418126090178654997034238923046320180008239051499490538421036244430389657609543220871622601848312332395555355812758453650812751650779322991406320835368022271567955630963981744522450178266909953191453192860426277757634233299308910808873088486615409217343470751281189670701718188980744852133602312807078578742518487429923088699783834193489412796969540792737023260804238965063062886656493672907540727939507037978464076527;
assign k3 = 1506'd249451153586847904964811286725161370143571293947219677900524009999253900587667899783359237764094121879966607070217086550289159163416107317632978859787150407791358079215752653065529229347009539469644878242563779410468386044030190551965974558003069521569385675851155169873444730578940738379571153338660041592616529376545020785682197847595605125610332701091477190740675966475331346435501040677175858692981081478349863476029841080244104079779347387600628355;
assign xo = 1506'd1166834498785274165882740778956565969045253728549738602599847879924360085539649388898405185185486720690454338894029385697558708490158429533023662699859451913087792442431648775012131670941338217306010447961839865076127582026944103049367477552558158300328503910891478772223197503338024587320433750019408976738770125318481870653333305634312799725972386027773574241887542793664878026780187760378733122398627276781066754263178210112265719209640365452406354828;
assign zo = 1506'd1396331324935382590778825339276267563026828108473684325109240786851362021089313714859780365535448442783041500434960909483279487331776481237256460709877882797417853329306815930754704327602710840640395023260234112244491886371492506737080921985849730146521562332872682701915005153911584790593871534987696096701419994081507516559046774869362328978183466281621171017360619955117263004577608446161756812793666190332127102801472249300390950504315518869873828062;

cryptoprocessor_wrapper_1506 UUT(clk,rst,get_output,data_en,ins_in,command_in,din_1,din_2,dout_1,dout_2);

always #1 clk = ~clk;

initial begin
    clk = 0; rst = 0; data_en = 0; ins_in = 0; get_output = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd0,7'd0,7'd0,7'd0};
    @(posedge clk);
    rst = 1;get_output = 0;
    @(posedge clk);
    rst = 0;
    @(posedge clk);
    //Load x in addr 0
    data_en = 1; ins_in = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd1,7'd0,7'd0,7'd0};
    din_1 = x;
    din_2 = 0;
    @(posedge clk);
    //Load z in addr 1
    data_en = 1; ins_in = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd1,7'd0,7'd0,7'd1};
    din_1 = z;
    din_2 = 0;
    @(posedge clk);
    //Load k1 in addr 2
    data_en = 1; ins_in = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd1,7'd0,7'd0,7'd2};
    din_1 = k1;
    din_2 = 0;
    @(posedge clk);
    //Load k2 in addr 3
    data_en = 1; ins_in = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd1,7'd0,7'd0,7'd3};
    din_1 = k2;
    din_2 = 0;
    @(posedge clk);
    //Load k3 in addr 4
    data_en = 1; ins_in = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd1,7'd0,7'd0,7'd4};
    din_1 = k3;
    din_2 = 0;
    @(posedge clk);
    
    //Start the operations
    //addr5 = addr0 + addr1 | t0 = x + z
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd3,7'd0,7'd1,7'd5};
    @(posedge clk);
    //addr6 = addr0 - addr1 | t1 = x - z
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd4,7'd0,7'd1,7'd6};
    @(posedge clk);
    //addr7 = addr5 * addr3 | x0 = t0 * K2
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd5,7'd3,7'd7};
    @(posedge clk);
    //addr8 = addr6 * addr4 | z0 = t1 * K3
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd6,7'd4,7'd8};
    @(posedge clk);
    //addr5 = addr5 * addr6 | t0 = t0 * t1
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd5,7'd6,7'd5};
    @(posedge clk);
    //addr5 = addr5 * addr2 | t0 = t0 * k1
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd5,7'd2,7'd5};
    @(posedge clk);
    //addr6 = addr7 + addr8 | t1 = xo + zo 
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd3,7'd7,7'd8,7'd6};
    @(posedge clk);
    //addr8 = addr7 - addr8 | zo = xo - zo   
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd4,7'd7,7'd8,7'd8};
    @(posedge clk);
    //addr6 = addr6 * addr6 | t1 = t1 * t1
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd6,7'd6,7'd6};
    @(posedge clk);
    //addr8 = addr8 * addr8 | zo = zo * zo 
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd8,7'd8,7'd8};
    @(posedge clk);
    //addr7 = addr5 + addr6 | xo = t0 + t1
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd3,7'd5,7'd6,7'd7};
    @(posedge clk);
    //addr5 = addr8 - addr5 | t0 = zo - t0
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd4,7'd8,7'd5,7'd5};
    @(posedge clk);
    //addr7 = addr7 * addr6 | xo = xo * t1
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd7,7'd6,7'd7};
    @(posedge clk);
    //addr8 = addr8 * addr5 | zo = zo * t0
    data_en = 0;ins_in = 1; din_1 = 0;din_2 = 0;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd5,7'd8,7'd5,7'd8};
    @(posedge clk);
    
    //Get output of addr = 7
    get_output = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd0,7'd7,7'd0,7'd0};
    @(posedge clk);
    if (xo != calculated) begin
        $display("TEST for 4_iso_c: FAILED.");
        $display("Failed TEST: output = 0x%x,0x%x | x->4_iso_c = 0x%x, calculated = 0x%x",dout_1,dout_2,xo,calculated);
        $display("Failed TEST: inputs: x,z = 0x%x,0x%x",x,z);
        $stop();
    end
    //Get output of addr = 8
    get_output = 1;
    {INS,rd_addr_1,rd_addr_2,wr_addr} = {3'd0,7'd8,7'd0,7'd0};
    @(posedge clk);
    if (zo != calculated) begin
        $display("TEST for 4_iso_c: FAILED.");
        $display("Failed TEST: output = 0x%x,0x%x | z->4_iso_c = 0x%x, calculated = 0x%x",dout_1,dout_2,zo,calculated);
        $display("Failed TEST: inputs: x,z = 0x%x,0x%x",x,z);
        $stop();
    end

    @(posedge clk);
    
    $display("4-iso-e correct");
    $finish();
end

endmodule
    