
module fa(
    input x,y,z,
    output c,s
);

assign {c,s} = x+y+z;

endmodule
    