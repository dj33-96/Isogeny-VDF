

module csa_tree_1506x3012(
    input [4536071:0] A, // lines are appended together
    output[3011:0] B_0,
    output[3011:0] B_1
);

wire [3024047:0] tree_1;
wire [2018039:0] tree_2;
wire [1346363:0] tree_3;
wire [897575:0] tree_4;
wire [599387:0] tree_5;
wire [400595:0] tree_6;
wire [268067:0] tree_7;
wire [180719:0] tree_8;
wire [120479:0] tree_9;
wire [81323:0] tree_10;
wire [54215:0] tree_11;
wire [36143:0] tree_12;
wire [24095:0] tree_13;
wire [18071:0] tree_14;
wire [12047:0] tree_15;
wire [9035:0] tree_16;
wire [6023:0] tree_17;
// layer-1
csa_3012 csau_3012_i0(A[3011:0],A[6023:3012],A[9035:6024],tree_1[3011:0],tree_1[6023:3012]);
csa_3012 csau_3012_i1(A[12047:9036],A[15059:12048],A[18071:15060],tree_1[9035:6024],tree_1[12047:9036]);
csa_3012 csau_3012_i2(A[21083:18072],A[24095:21084],A[27107:24096],tree_1[15059:12048],tree_1[18071:15060]);
csa_3012 csau_3012_i3(A[30119:27108],A[33131:30120],A[36143:33132],tree_1[21083:18072],tree_1[24095:21084]);
csa_3012 csau_3012_i4(A[39155:36144],A[42167:39156],A[45179:42168],tree_1[27107:24096],tree_1[30119:27108]);
csa_3012 csau_3012_i5(A[48191:45180],A[51203:48192],A[54215:51204],tree_1[33131:30120],tree_1[36143:33132]);
csa_3012 csau_3012_i6(A[57227:54216],A[60239:57228],A[63251:60240],tree_1[39155:36144],tree_1[42167:39156]);
csa_3012 csau_3012_i7(A[66263:63252],A[69275:66264],A[72287:69276],tree_1[45179:42168],tree_1[48191:45180]);
csa_3012 csau_3012_i8(A[75299:72288],A[78311:75300],A[81323:78312],tree_1[51203:48192],tree_1[54215:51204]);
csa_3012 csau_3012_i9(A[84335:81324],A[87347:84336],A[90359:87348],tree_1[57227:54216],tree_1[60239:57228]);
csa_3012 csau_3012_i10(A[93371:90360],A[96383:93372],A[99395:96384],tree_1[63251:60240],tree_1[66263:63252]);
csa_3012 csau_3012_i11(A[102407:99396],A[105419:102408],A[108431:105420],tree_1[69275:66264],tree_1[72287:69276]);
csa_3012 csau_3012_i12(A[111443:108432],A[114455:111444],A[117467:114456],tree_1[75299:72288],tree_1[78311:75300]);
csa_3012 csau_3012_i13(A[120479:117468],A[123491:120480],A[126503:123492],tree_1[81323:78312],tree_1[84335:81324]);
csa_3012 csau_3012_i14(A[129515:126504],A[132527:129516],A[135539:132528],tree_1[87347:84336],tree_1[90359:87348]);
csa_3012 csau_3012_i15(A[138551:135540],A[141563:138552],A[144575:141564],tree_1[93371:90360],tree_1[96383:93372]);
csa_3012 csau_3012_i16(A[147587:144576],A[150599:147588],A[153611:150600],tree_1[99395:96384],tree_1[102407:99396]);
csa_3012 csau_3012_i17(A[156623:153612],A[159635:156624],A[162647:159636],tree_1[105419:102408],tree_1[108431:105420]);
csa_3012 csau_3012_i18(A[165659:162648],A[168671:165660],A[171683:168672],tree_1[111443:108432],tree_1[114455:111444]);
csa_3012 csau_3012_i19(A[174695:171684],A[177707:174696],A[180719:177708],tree_1[117467:114456],tree_1[120479:117468]);
csa_3012 csau_3012_i20(A[183731:180720],A[186743:183732],A[189755:186744],tree_1[123491:120480],tree_1[126503:123492]);
csa_3012 csau_3012_i21(A[192767:189756],A[195779:192768],A[198791:195780],tree_1[129515:126504],tree_1[132527:129516]);
csa_3012 csau_3012_i22(A[201803:198792],A[204815:201804],A[207827:204816],tree_1[135539:132528],tree_1[138551:135540]);
csa_3012 csau_3012_i23(A[210839:207828],A[213851:210840],A[216863:213852],tree_1[141563:138552],tree_1[144575:141564]);
csa_3012 csau_3012_i24(A[219875:216864],A[222887:219876],A[225899:222888],tree_1[147587:144576],tree_1[150599:147588]);
csa_3012 csau_3012_i25(A[228911:225900],A[231923:228912],A[234935:231924],tree_1[153611:150600],tree_1[156623:153612]);
csa_3012 csau_3012_i26(A[237947:234936],A[240959:237948],A[243971:240960],tree_1[159635:156624],tree_1[162647:159636]);
csa_3012 csau_3012_i27(A[246983:243972],A[249995:246984],A[253007:249996],tree_1[165659:162648],tree_1[168671:165660]);
csa_3012 csau_3012_i28(A[256019:253008],A[259031:256020],A[262043:259032],tree_1[171683:168672],tree_1[174695:171684]);
csa_3012 csau_3012_i29(A[265055:262044],A[268067:265056],A[271079:268068],tree_1[177707:174696],tree_1[180719:177708]);
csa_3012 csau_3012_i30(A[274091:271080],A[277103:274092],A[280115:277104],tree_1[183731:180720],tree_1[186743:183732]);
csa_3012 csau_3012_i31(A[283127:280116],A[286139:283128],A[289151:286140],tree_1[189755:186744],tree_1[192767:189756]);
csa_3012 csau_3012_i32(A[292163:289152],A[295175:292164],A[298187:295176],tree_1[195779:192768],tree_1[198791:195780]);
csa_3012 csau_3012_i33(A[301199:298188],A[304211:301200],A[307223:304212],tree_1[201803:198792],tree_1[204815:201804]);
csa_3012 csau_3012_i34(A[310235:307224],A[313247:310236],A[316259:313248],tree_1[207827:204816],tree_1[210839:207828]);
csa_3012 csau_3012_i35(A[319271:316260],A[322283:319272],A[325295:322284],tree_1[213851:210840],tree_1[216863:213852]);
csa_3012 csau_3012_i36(A[328307:325296],A[331319:328308],A[334331:331320],tree_1[219875:216864],tree_1[222887:219876]);
csa_3012 csau_3012_i37(A[337343:334332],A[340355:337344],A[343367:340356],tree_1[225899:222888],tree_1[228911:225900]);
csa_3012 csau_3012_i38(A[346379:343368],A[349391:346380],A[352403:349392],tree_1[231923:228912],tree_1[234935:231924]);
csa_3012 csau_3012_i39(A[355415:352404],A[358427:355416],A[361439:358428],tree_1[237947:234936],tree_1[240959:237948]);
csa_3012 csau_3012_i40(A[364451:361440],A[367463:364452],A[370475:367464],tree_1[243971:240960],tree_1[246983:243972]);
csa_3012 csau_3012_i41(A[373487:370476],A[376499:373488],A[379511:376500],tree_1[249995:246984],tree_1[253007:249996]);
csa_3012 csau_3012_i42(A[382523:379512],A[385535:382524],A[388547:385536],tree_1[256019:253008],tree_1[259031:256020]);
csa_3012 csau_3012_i43(A[391559:388548],A[394571:391560],A[397583:394572],tree_1[262043:259032],tree_1[265055:262044]);
csa_3012 csau_3012_i44(A[400595:397584],A[403607:400596],A[406619:403608],tree_1[268067:265056],tree_1[271079:268068]);
csa_3012 csau_3012_i45(A[409631:406620],A[412643:409632],A[415655:412644],tree_1[274091:271080],tree_1[277103:274092]);
csa_3012 csau_3012_i46(A[418667:415656],A[421679:418668],A[424691:421680],tree_1[280115:277104],tree_1[283127:280116]);
csa_3012 csau_3012_i47(A[427703:424692],A[430715:427704],A[433727:430716],tree_1[286139:283128],tree_1[289151:286140]);
csa_3012 csau_3012_i48(A[436739:433728],A[439751:436740],A[442763:439752],tree_1[292163:289152],tree_1[295175:292164]);
csa_3012 csau_3012_i49(A[445775:442764],A[448787:445776],A[451799:448788],tree_1[298187:295176],tree_1[301199:298188]);
csa_3012 csau_3012_i50(A[454811:451800],A[457823:454812],A[460835:457824],tree_1[304211:301200],tree_1[307223:304212]);
csa_3012 csau_3012_i51(A[463847:460836],A[466859:463848],A[469871:466860],tree_1[310235:307224],tree_1[313247:310236]);
csa_3012 csau_3012_i52(A[472883:469872],A[475895:472884],A[478907:475896],tree_1[316259:313248],tree_1[319271:316260]);
csa_3012 csau_3012_i53(A[481919:478908],A[484931:481920],A[487943:484932],tree_1[322283:319272],tree_1[325295:322284]);
csa_3012 csau_3012_i54(A[490955:487944],A[493967:490956],A[496979:493968],tree_1[328307:325296],tree_1[331319:328308]);
csa_3012 csau_3012_i55(A[499991:496980],A[503003:499992],A[506015:503004],tree_1[334331:331320],tree_1[337343:334332]);
csa_3012 csau_3012_i56(A[509027:506016],A[512039:509028],A[515051:512040],tree_1[340355:337344],tree_1[343367:340356]);
csa_3012 csau_3012_i57(A[518063:515052],A[521075:518064],A[524087:521076],tree_1[346379:343368],tree_1[349391:346380]);
csa_3012 csau_3012_i58(A[527099:524088],A[530111:527100],A[533123:530112],tree_1[352403:349392],tree_1[355415:352404]);
csa_3012 csau_3012_i59(A[536135:533124],A[539147:536136],A[542159:539148],tree_1[358427:355416],tree_1[361439:358428]);
csa_3012 csau_3012_i60(A[545171:542160],A[548183:545172],A[551195:548184],tree_1[364451:361440],tree_1[367463:364452]);
csa_3012 csau_3012_i61(A[554207:551196],A[557219:554208],A[560231:557220],tree_1[370475:367464],tree_1[373487:370476]);
csa_3012 csau_3012_i62(A[563243:560232],A[566255:563244],A[569267:566256],tree_1[376499:373488],tree_1[379511:376500]);
csa_3012 csau_3012_i63(A[572279:569268],A[575291:572280],A[578303:575292],tree_1[382523:379512],tree_1[385535:382524]);
csa_3012 csau_3012_i64(A[581315:578304],A[584327:581316],A[587339:584328],tree_1[388547:385536],tree_1[391559:388548]);
csa_3012 csau_3012_i65(A[590351:587340],A[593363:590352],A[596375:593364],tree_1[394571:391560],tree_1[397583:394572]);
csa_3012 csau_3012_i66(A[599387:596376],A[602399:599388],A[605411:602400],tree_1[400595:397584],tree_1[403607:400596]);
csa_3012 csau_3012_i67(A[608423:605412],A[611435:608424],A[614447:611436],tree_1[406619:403608],tree_1[409631:406620]);
csa_3012 csau_3012_i68(A[617459:614448],A[620471:617460],A[623483:620472],tree_1[412643:409632],tree_1[415655:412644]);
csa_3012 csau_3012_i69(A[626495:623484],A[629507:626496],A[632519:629508],tree_1[418667:415656],tree_1[421679:418668]);
csa_3012 csau_3012_i70(A[635531:632520],A[638543:635532],A[641555:638544],tree_1[424691:421680],tree_1[427703:424692]);
csa_3012 csau_3012_i71(A[644567:641556],A[647579:644568],A[650591:647580],tree_1[430715:427704],tree_1[433727:430716]);
csa_3012 csau_3012_i72(A[653603:650592],A[656615:653604],A[659627:656616],tree_1[436739:433728],tree_1[439751:436740]);
csa_3012 csau_3012_i73(A[662639:659628],A[665651:662640],A[668663:665652],tree_1[442763:439752],tree_1[445775:442764]);
csa_3012 csau_3012_i74(A[671675:668664],A[674687:671676],A[677699:674688],tree_1[448787:445776],tree_1[451799:448788]);
csa_3012 csau_3012_i75(A[680711:677700],A[683723:680712],A[686735:683724],tree_1[454811:451800],tree_1[457823:454812]);
csa_3012 csau_3012_i76(A[689747:686736],A[692759:689748],A[695771:692760],tree_1[460835:457824],tree_1[463847:460836]);
csa_3012 csau_3012_i77(A[698783:695772],A[701795:698784],A[704807:701796],tree_1[466859:463848],tree_1[469871:466860]);
csa_3012 csau_3012_i78(A[707819:704808],A[710831:707820],A[713843:710832],tree_1[472883:469872],tree_1[475895:472884]);
csa_3012 csau_3012_i79(A[716855:713844],A[719867:716856],A[722879:719868],tree_1[478907:475896],tree_1[481919:478908]);
csa_3012 csau_3012_i80(A[725891:722880],A[728903:725892],A[731915:728904],tree_1[484931:481920],tree_1[487943:484932]);
csa_3012 csau_3012_i81(A[734927:731916],A[737939:734928],A[740951:737940],tree_1[490955:487944],tree_1[493967:490956]);
csa_3012 csau_3012_i82(A[743963:740952],A[746975:743964],A[749987:746976],tree_1[496979:493968],tree_1[499991:496980]);
csa_3012 csau_3012_i83(A[752999:749988],A[756011:753000],A[759023:756012],tree_1[503003:499992],tree_1[506015:503004]);
csa_3012 csau_3012_i84(A[762035:759024],A[765047:762036],A[768059:765048],tree_1[509027:506016],tree_1[512039:509028]);
csa_3012 csau_3012_i85(A[771071:768060],A[774083:771072],A[777095:774084],tree_1[515051:512040],tree_1[518063:515052]);
csa_3012 csau_3012_i86(A[780107:777096],A[783119:780108],A[786131:783120],tree_1[521075:518064],tree_1[524087:521076]);
csa_3012 csau_3012_i87(A[789143:786132],A[792155:789144],A[795167:792156],tree_1[527099:524088],tree_1[530111:527100]);
csa_3012 csau_3012_i88(A[798179:795168],A[801191:798180],A[804203:801192],tree_1[533123:530112],tree_1[536135:533124]);
csa_3012 csau_3012_i89(A[807215:804204],A[810227:807216],A[813239:810228],tree_1[539147:536136],tree_1[542159:539148]);
csa_3012 csau_3012_i90(A[816251:813240],A[819263:816252],A[822275:819264],tree_1[545171:542160],tree_1[548183:545172]);
csa_3012 csau_3012_i91(A[825287:822276],A[828299:825288],A[831311:828300],tree_1[551195:548184],tree_1[554207:551196]);
csa_3012 csau_3012_i92(A[834323:831312],A[837335:834324],A[840347:837336],tree_1[557219:554208],tree_1[560231:557220]);
csa_3012 csau_3012_i93(A[843359:840348],A[846371:843360],A[849383:846372],tree_1[563243:560232],tree_1[566255:563244]);
csa_3012 csau_3012_i94(A[852395:849384],A[855407:852396],A[858419:855408],tree_1[569267:566256],tree_1[572279:569268]);
csa_3012 csau_3012_i95(A[861431:858420],A[864443:861432],A[867455:864444],tree_1[575291:572280],tree_1[578303:575292]);
csa_3012 csau_3012_i96(A[870467:867456],A[873479:870468],A[876491:873480],tree_1[581315:578304],tree_1[584327:581316]);
csa_3012 csau_3012_i97(A[879503:876492],A[882515:879504],A[885527:882516],tree_1[587339:584328],tree_1[590351:587340]);
csa_3012 csau_3012_i98(A[888539:885528],A[891551:888540],A[894563:891552],tree_1[593363:590352],tree_1[596375:593364]);
csa_3012 csau_3012_i99(A[897575:894564],A[900587:897576],A[903599:900588],tree_1[599387:596376],tree_1[602399:599388]);
csa_3012 csau_3012_i100(A[906611:903600],A[909623:906612],A[912635:909624],tree_1[605411:602400],tree_1[608423:605412]);
csa_3012 csau_3012_i101(A[915647:912636],A[918659:915648],A[921671:918660],tree_1[611435:608424],tree_1[614447:611436]);
csa_3012 csau_3012_i102(A[924683:921672],A[927695:924684],A[930707:927696],tree_1[617459:614448],tree_1[620471:617460]);
csa_3012 csau_3012_i103(A[933719:930708],A[936731:933720],A[939743:936732],tree_1[623483:620472],tree_1[626495:623484]);
csa_3012 csau_3012_i104(A[942755:939744],A[945767:942756],A[948779:945768],tree_1[629507:626496],tree_1[632519:629508]);
csa_3012 csau_3012_i105(A[951791:948780],A[954803:951792],A[957815:954804],tree_1[635531:632520],tree_1[638543:635532]);
csa_3012 csau_3012_i106(A[960827:957816],A[963839:960828],A[966851:963840],tree_1[641555:638544],tree_1[644567:641556]);
csa_3012 csau_3012_i107(A[969863:966852],A[972875:969864],A[975887:972876],tree_1[647579:644568],tree_1[650591:647580]);
csa_3012 csau_3012_i108(A[978899:975888],A[981911:978900],A[984923:981912],tree_1[653603:650592],tree_1[656615:653604]);
csa_3012 csau_3012_i109(A[987935:984924],A[990947:987936],A[993959:990948],tree_1[659627:656616],tree_1[662639:659628]);
csa_3012 csau_3012_i110(A[996971:993960],A[999983:996972],A[1002995:999984],tree_1[665651:662640],tree_1[668663:665652]);
csa_3012 csau_3012_i111(A[1006007:1002996],A[1009019:1006008],A[1012031:1009020],tree_1[671675:668664],tree_1[674687:671676]);
csa_3012 csau_3012_i112(A[1015043:1012032],A[1018055:1015044],A[1021067:1018056],tree_1[677699:674688],tree_1[680711:677700]);
csa_3012 csau_3012_i113(A[1024079:1021068],A[1027091:1024080],A[1030103:1027092],tree_1[683723:680712],tree_1[686735:683724]);
csa_3012 csau_3012_i114(A[1033115:1030104],A[1036127:1033116],A[1039139:1036128],tree_1[689747:686736],tree_1[692759:689748]);
csa_3012 csau_3012_i115(A[1042151:1039140],A[1045163:1042152],A[1048175:1045164],tree_1[695771:692760],tree_1[698783:695772]);
csa_3012 csau_3012_i116(A[1051187:1048176],A[1054199:1051188],A[1057211:1054200],tree_1[701795:698784],tree_1[704807:701796]);
csa_3012 csau_3012_i117(A[1060223:1057212],A[1063235:1060224],A[1066247:1063236],tree_1[707819:704808],tree_1[710831:707820]);
csa_3012 csau_3012_i118(A[1069259:1066248],A[1072271:1069260],A[1075283:1072272],tree_1[713843:710832],tree_1[716855:713844]);
csa_3012 csau_3012_i119(A[1078295:1075284],A[1081307:1078296],A[1084319:1081308],tree_1[719867:716856],tree_1[722879:719868]);
csa_3012 csau_3012_i120(A[1087331:1084320],A[1090343:1087332],A[1093355:1090344],tree_1[725891:722880],tree_1[728903:725892]);
csa_3012 csau_3012_i121(A[1096367:1093356],A[1099379:1096368],A[1102391:1099380],tree_1[731915:728904],tree_1[734927:731916]);
csa_3012 csau_3012_i122(A[1105403:1102392],A[1108415:1105404],A[1111427:1108416],tree_1[737939:734928],tree_1[740951:737940]);
csa_3012 csau_3012_i123(A[1114439:1111428],A[1117451:1114440],A[1120463:1117452],tree_1[743963:740952],tree_1[746975:743964]);
csa_3012 csau_3012_i124(A[1123475:1120464],A[1126487:1123476],A[1129499:1126488],tree_1[749987:746976],tree_1[752999:749988]);
csa_3012 csau_3012_i125(A[1132511:1129500],A[1135523:1132512],A[1138535:1135524],tree_1[756011:753000],tree_1[759023:756012]);
csa_3012 csau_3012_i126(A[1141547:1138536],A[1144559:1141548],A[1147571:1144560],tree_1[762035:759024],tree_1[765047:762036]);
csa_3012 csau_3012_i127(A[1150583:1147572],A[1153595:1150584],A[1156607:1153596],tree_1[768059:765048],tree_1[771071:768060]);
csa_3012 csau_3012_i128(A[1159619:1156608],A[1162631:1159620],A[1165643:1162632],tree_1[774083:771072],tree_1[777095:774084]);
csa_3012 csau_3012_i129(A[1168655:1165644],A[1171667:1168656],A[1174679:1171668],tree_1[780107:777096],tree_1[783119:780108]);
csa_3012 csau_3012_i130(A[1177691:1174680],A[1180703:1177692],A[1183715:1180704],tree_1[786131:783120],tree_1[789143:786132]);
csa_3012 csau_3012_i131(A[1186727:1183716],A[1189739:1186728],A[1192751:1189740],tree_1[792155:789144],tree_1[795167:792156]);
csa_3012 csau_3012_i132(A[1195763:1192752],A[1198775:1195764],A[1201787:1198776],tree_1[798179:795168],tree_1[801191:798180]);
csa_3012 csau_3012_i133(A[1204799:1201788],A[1207811:1204800],A[1210823:1207812],tree_1[804203:801192],tree_1[807215:804204]);
csa_3012 csau_3012_i134(A[1213835:1210824],A[1216847:1213836],A[1219859:1216848],tree_1[810227:807216],tree_1[813239:810228]);
csa_3012 csau_3012_i135(A[1222871:1219860],A[1225883:1222872],A[1228895:1225884],tree_1[816251:813240],tree_1[819263:816252]);
csa_3012 csau_3012_i136(A[1231907:1228896],A[1234919:1231908],A[1237931:1234920],tree_1[822275:819264],tree_1[825287:822276]);
csa_3012 csau_3012_i137(A[1240943:1237932],A[1243955:1240944],A[1246967:1243956],tree_1[828299:825288],tree_1[831311:828300]);
csa_3012 csau_3012_i138(A[1249979:1246968],A[1252991:1249980],A[1256003:1252992],tree_1[834323:831312],tree_1[837335:834324]);
csa_3012 csau_3012_i139(A[1259015:1256004],A[1262027:1259016],A[1265039:1262028],tree_1[840347:837336],tree_1[843359:840348]);
csa_3012 csau_3012_i140(A[1268051:1265040],A[1271063:1268052],A[1274075:1271064],tree_1[846371:843360],tree_1[849383:846372]);
csa_3012 csau_3012_i141(A[1277087:1274076],A[1280099:1277088],A[1283111:1280100],tree_1[852395:849384],tree_1[855407:852396]);
csa_3012 csau_3012_i142(A[1286123:1283112],A[1289135:1286124],A[1292147:1289136],tree_1[858419:855408],tree_1[861431:858420]);
csa_3012 csau_3012_i143(A[1295159:1292148],A[1298171:1295160],A[1301183:1298172],tree_1[864443:861432],tree_1[867455:864444]);
csa_3012 csau_3012_i144(A[1304195:1301184],A[1307207:1304196],A[1310219:1307208],tree_1[870467:867456],tree_1[873479:870468]);
csa_3012 csau_3012_i145(A[1313231:1310220],A[1316243:1313232],A[1319255:1316244],tree_1[876491:873480],tree_1[879503:876492]);
csa_3012 csau_3012_i146(A[1322267:1319256],A[1325279:1322268],A[1328291:1325280],tree_1[882515:879504],tree_1[885527:882516]);
csa_3012 csau_3012_i147(A[1331303:1328292],A[1334315:1331304],A[1337327:1334316],tree_1[888539:885528],tree_1[891551:888540]);
csa_3012 csau_3012_i148(A[1340339:1337328],A[1343351:1340340],A[1346363:1343352],tree_1[894563:891552],tree_1[897575:894564]);
csa_3012 csau_3012_i149(A[1349375:1346364],A[1352387:1349376],A[1355399:1352388],tree_1[900587:897576],tree_1[903599:900588]);
csa_3012 csau_3012_i150(A[1358411:1355400],A[1361423:1358412],A[1364435:1361424],tree_1[906611:903600],tree_1[909623:906612]);
csa_3012 csau_3012_i151(A[1367447:1364436],A[1370459:1367448],A[1373471:1370460],tree_1[912635:909624],tree_1[915647:912636]);
csa_3012 csau_3012_i152(A[1376483:1373472],A[1379495:1376484],A[1382507:1379496],tree_1[918659:915648],tree_1[921671:918660]);
csa_3012 csau_3012_i153(A[1385519:1382508],A[1388531:1385520],A[1391543:1388532],tree_1[924683:921672],tree_1[927695:924684]);
csa_3012 csau_3012_i154(A[1394555:1391544],A[1397567:1394556],A[1400579:1397568],tree_1[930707:927696],tree_1[933719:930708]);
csa_3012 csau_3012_i155(A[1403591:1400580],A[1406603:1403592],A[1409615:1406604],tree_1[936731:933720],tree_1[939743:936732]);
csa_3012 csau_3012_i156(A[1412627:1409616],A[1415639:1412628],A[1418651:1415640],tree_1[942755:939744],tree_1[945767:942756]);
csa_3012 csau_3012_i157(A[1421663:1418652],A[1424675:1421664],A[1427687:1424676],tree_1[948779:945768],tree_1[951791:948780]);
csa_3012 csau_3012_i158(A[1430699:1427688],A[1433711:1430700],A[1436723:1433712],tree_1[954803:951792],tree_1[957815:954804]);
csa_3012 csau_3012_i159(A[1439735:1436724],A[1442747:1439736],A[1445759:1442748],tree_1[960827:957816],tree_1[963839:960828]);
csa_3012 csau_3012_i160(A[1448771:1445760],A[1451783:1448772],A[1454795:1451784],tree_1[966851:963840],tree_1[969863:966852]);
csa_3012 csau_3012_i161(A[1457807:1454796],A[1460819:1457808],A[1463831:1460820],tree_1[972875:969864],tree_1[975887:972876]);
csa_3012 csau_3012_i162(A[1466843:1463832],A[1469855:1466844],A[1472867:1469856],tree_1[978899:975888],tree_1[981911:978900]);
csa_3012 csau_3012_i163(A[1475879:1472868],A[1478891:1475880],A[1481903:1478892],tree_1[984923:981912],tree_1[987935:984924]);
csa_3012 csau_3012_i164(A[1484915:1481904],A[1487927:1484916],A[1490939:1487928],tree_1[990947:987936],tree_1[993959:990948]);
csa_3012 csau_3012_i165(A[1493951:1490940],A[1496963:1493952],A[1499975:1496964],tree_1[996971:993960],tree_1[999983:996972]);
csa_3012 csau_3012_i166(A[1502987:1499976],A[1505999:1502988],A[1509011:1506000],tree_1[1002995:999984],tree_1[1006007:1002996]);
csa_3012 csau_3012_i167(A[1512023:1509012],A[1515035:1512024],A[1518047:1515036],tree_1[1009019:1006008],tree_1[1012031:1009020]);
csa_3012 csau_3012_i168(A[1521059:1518048],A[1524071:1521060],A[1527083:1524072],tree_1[1015043:1012032],tree_1[1018055:1015044]);
csa_3012 csau_3012_i169(A[1530095:1527084],A[1533107:1530096],A[1536119:1533108],tree_1[1021067:1018056],tree_1[1024079:1021068]);
csa_3012 csau_3012_i170(A[1539131:1536120],A[1542143:1539132],A[1545155:1542144],tree_1[1027091:1024080],tree_1[1030103:1027092]);
csa_3012 csau_3012_i171(A[1548167:1545156],A[1551179:1548168],A[1554191:1551180],tree_1[1033115:1030104],tree_1[1036127:1033116]);
csa_3012 csau_3012_i172(A[1557203:1554192],A[1560215:1557204],A[1563227:1560216],tree_1[1039139:1036128],tree_1[1042151:1039140]);
csa_3012 csau_3012_i173(A[1566239:1563228],A[1569251:1566240],A[1572263:1569252],tree_1[1045163:1042152],tree_1[1048175:1045164]);
csa_3012 csau_3012_i174(A[1575275:1572264],A[1578287:1575276],A[1581299:1578288],tree_1[1051187:1048176],tree_1[1054199:1051188]);
csa_3012 csau_3012_i175(A[1584311:1581300],A[1587323:1584312],A[1590335:1587324],tree_1[1057211:1054200],tree_1[1060223:1057212]);
csa_3012 csau_3012_i176(A[1593347:1590336],A[1596359:1593348],A[1599371:1596360],tree_1[1063235:1060224],tree_1[1066247:1063236]);
csa_3012 csau_3012_i177(A[1602383:1599372],A[1605395:1602384],A[1608407:1605396],tree_1[1069259:1066248],tree_1[1072271:1069260]);
csa_3012 csau_3012_i178(A[1611419:1608408],A[1614431:1611420],A[1617443:1614432],tree_1[1075283:1072272],tree_1[1078295:1075284]);
csa_3012 csau_3012_i179(A[1620455:1617444],A[1623467:1620456],A[1626479:1623468],tree_1[1081307:1078296],tree_1[1084319:1081308]);
csa_3012 csau_3012_i180(A[1629491:1626480],A[1632503:1629492],A[1635515:1632504],tree_1[1087331:1084320],tree_1[1090343:1087332]);
csa_3012 csau_3012_i181(A[1638527:1635516],A[1641539:1638528],A[1644551:1641540],tree_1[1093355:1090344],tree_1[1096367:1093356]);
csa_3012 csau_3012_i182(A[1647563:1644552],A[1650575:1647564],A[1653587:1650576],tree_1[1099379:1096368],tree_1[1102391:1099380]);
csa_3012 csau_3012_i183(A[1656599:1653588],A[1659611:1656600],A[1662623:1659612],tree_1[1105403:1102392],tree_1[1108415:1105404]);
csa_3012 csau_3012_i184(A[1665635:1662624],A[1668647:1665636],A[1671659:1668648],tree_1[1111427:1108416],tree_1[1114439:1111428]);
csa_3012 csau_3012_i185(A[1674671:1671660],A[1677683:1674672],A[1680695:1677684],tree_1[1117451:1114440],tree_1[1120463:1117452]);
csa_3012 csau_3012_i186(A[1683707:1680696],A[1686719:1683708],A[1689731:1686720],tree_1[1123475:1120464],tree_1[1126487:1123476]);
csa_3012 csau_3012_i187(A[1692743:1689732],A[1695755:1692744],A[1698767:1695756],tree_1[1129499:1126488],tree_1[1132511:1129500]);
csa_3012 csau_3012_i188(A[1701779:1698768],A[1704791:1701780],A[1707803:1704792],tree_1[1135523:1132512],tree_1[1138535:1135524]);
csa_3012 csau_3012_i189(A[1710815:1707804],A[1713827:1710816],A[1716839:1713828],tree_1[1141547:1138536],tree_1[1144559:1141548]);
csa_3012 csau_3012_i190(A[1719851:1716840],A[1722863:1719852],A[1725875:1722864],tree_1[1147571:1144560],tree_1[1150583:1147572]);
csa_3012 csau_3012_i191(A[1728887:1725876],A[1731899:1728888],A[1734911:1731900],tree_1[1153595:1150584],tree_1[1156607:1153596]);
csa_3012 csau_3012_i192(A[1737923:1734912],A[1740935:1737924],A[1743947:1740936],tree_1[1159619:1156608],tree_1[1162631:1159620]);
csa_3012 csau_3012_i193(A[1746959:1743948],A[1749971:1746960],A[1752983:1749972],tree_1[1165643:1162632],tree_1[1168655:1165644]);
csa_3012 csau_3012_i194(A[1755995:1752984],A[1759007:1755996],A[1762019:1759008],tree_1[1171667:1168656],tree_1[1174679:1171668]);
csa_3012 csau_3012_i195(A[1765031:1762020],A[1768043:1765032],A[1771055:1768044],tree_1[1177691:1174680],tree_1[1180703:1177692]);
csa_3012 csau_3012_i196(A[1774067:1771056],A[1777079:1774068],A[1780091:1777080],tree_1[1183715:1180704],tree_1[1186727:1183716]);
csa_3012 csau_3012_i197(A[1783103:1780092],A[1786115:1783104],A[1789127:1786116],tree_1[1189739:1186728],tree_1[1192751:1189740]);
csa_3012 csau_3012_i198(A[1792139:1789128],A[1795151:1792140],A[1798163:1795152],tree_1[1195763:1192752],tree_1[1198775:1195764]);
csa_3012 csau_3012_i199(A[1801175:1798164],A[1804187:1801176],A[1807199:1804188],tree_1[1201787:1198776],tree_1[1204799:1201788]);
csa_3012 csau_3012_i200(A[1810211:1807200],A[1813223:1810212],A[1816235:1813224],tree_1[1207811:1204800],tree_1[1210823:1207812]);
csa_3012 csau_3012_i201(A[1819247:1816236],A[1822259:1819248],A[1825271:1822260],tree_1[1213835:1210824],tree_1[1216847:1213836]);
csa_3012 csau_3012_i202(A[1828283:1825272],A[1831295:1828284],A[1834307:1831296],tree_1[1219859:1216848],tree_1[1222871:1219860]);
csa_3012 csau_3012_i203(A[1837319:1834308],A[1840331:1837320],A[1843343:1840332],tree_1[1225883:1222872],tree_1[1228895:1225884]);
csa_3012 csau_3012_i204(A[1846355:1843344],A[1849367:1846356],A[1852379:1849368],tree_1[1231907:1228896],tree_1[1234919:1231908]);
csa_3012 csau_3012_i205(A[1855391:1852380],A[1858403:1855392],A[1861415:1858404],tree_1[1237931:1234920],tree_1[1240943:1237932]);
csa_3012 csau_3012_i206(A[1864427:1861416],A[1867439:1864428],A[1870451:1867440],tree_1[1243955:1240944],tree_1[1246967:1243956]);
csa_3012 csau_3012_i207(A[1873463:1870452],A[1876475:1873464],A[1879487:1876476],tree_1[1249979:1246968],tree_1[1252991:1249980]);
csa_3012 csau_3012_i208(A[1882499:1879488],A[1885511:1882500],A[1888523:1885512],tree_1[1256003:1252992],tree_1[1259015:1256004]);
csa_3012 csau_3012_i209(A[1891535:1888524],A[1894547:1891536],A[1897559:1894548],tree_1[1262027:1259016],tree_1[1265039:1262028]);
csa_3012 csau_3012_i210(A[1900571:1897560],A[1903583:1900572],A[1906595:1903584],tree_1[1268051:1265040],tree_1[1271063:1268052]);
csa_3012 csau_3012_i211(A[1909607:1906596],A[1912619:1909608],A[1915631:1912620],tree_1[1274075:1271064],tree_1[1277087:1274076]);
csa_3012 csau_3012_i212(A[1918643:1915632],A[1921655:1918644],A[1924667:1921656],tree_1[1280099:1277088],tree_1[1283111:1280100]);
csa_3012 csau_3012_i213(A[1927679:1924668],A[1930691:1927680],A[1933703:1930692],tree_1[1286123:1283112],tree_1[1289135:1286124]);
csa_3012 csau_3012_i214(A[1936715:1933704],A[1939727:1936716],A[1942739:1939728],tree_1[1292147:1289136],tree_1[1295159:1292148]);
csa_3012 csau_3012_i215(A[1945751:1942740],A[1948763:1945752],A[1951775:1948764],tree_1[1298171:1295160],tree_1[1301183:1298172]);
csa_3012 csau_3012_i216(A[1954787:1951776],A[1957799:1954788],A[1960811:1957800],tree_1[1304195:1301184],tree_1[1307207:1304196]);
csa_3012 csau_3012_i217(A[1963823:1960812],A[1966835:1963824],A[1969847:1966836],tree_1[1310219:1307208],tree_1[1313231:1310220]);
csa_3012 csau_3012_i218(A[1972859:1969848],A[1975871:1972860],A[1978883:1975872],tree_1[1316243:1313232],tree_1[1319255:1316244]);
csa_3012 csau_3012_i219(A[1981895:1978884],A[1984907:1981896],A[1987919:1984908],tree_1[1322267:1319256],tree_1[1325279:1322268]);
csa_3012 csau_3012_i220(A[1990931:1987920],A[1993943:1990932],A[1996955:1993944],tree_1[1328291:1325280],tree_1[1331303:1328292]);
csa_3012 csau_3012_i221(A[1999967:1996956],A[2002979:1999968],A[2005991:2002980],tree_1[1334315:1331304],tree_1[1337327:1334316]);
csa_3012 csau_3012_i222(A[2009003:2005992],A[2012015:2009004],A[2015027:2012016],tree_1[1340339:1337328],tree_1[1343351:1340340]);
csa_3012 csau_3012_i223(A[2018039:2015028],A[2021051:2018040],A[2024063:2021052],tree_1[1346363:1343352],tree_1[1349375:1346364]);
csa_3012 csau_3012_i224(A[2027075:2024064],A[2030087:2027076],A[2033099:2030088],tree_1[1352387:1349376],tree_1[1355399:1352388]);
csa_3012 csau_3012_i225(A[2036111:2033100],A[2039123:2036112],A[2042135:2039124],tree_1[1358411:1355400],tree_1[1361423:1358412]);
csa_3012 csau_3012_i226(A[2045147:2042136],A[2048159:2045148],A[2051171:2048160],tree_1[1364435:1361424],tree_1[1367447:1364436]);
csa_3012 csau_3012_i227(A[2054183:2051172],A[2057195:2054184],A[2060207:2057196],tree_1[1370459:1367448],tree_1[1373471:1370460]);
csa_3012 csau_3012_i228(A[2063219:2060208],A[2066231:2063220],A[2069243:2066232],tree_1[1376483:1373472],tree_1[1379495:1376484]);
csa_3012 csau_3012_i229(A[2072255:2069244],A[2075267:2072256],A[2078279:2075268],tree_1[1382507:1379496],tree_1[1385519:1382508]);
csa_3012 csau_3012_i230(A[2081291:2078280],A[2084303:2081292],A[2087315:2084304],tree_1[1388531:1385520],tree_1[1391543:1388532]);
csa_3012 csau_3012_i231(A[2090327:2087316],A[2093339:2090328],A[2096351:2093340],tree_1[1394555:1391544],tree_1[1397567:1394556]);
csa_3012 csau_3012_i232(A[2099363:2096352],A[2102375:2099364],A[2105387:2102376],tree_1[1400579:1397568],tree_1[1403591:1400580]);
csa_3012 csau_3012_i233(A[2108399:2105388],A[2111411:2108400],A[2114423:2111412],tree_1[1406603:1403592],tree_1[1409615:1406604]);
csa_3012 csau_3012_i234(A[2117435:2114424],A[2120447:2117436],A[2123459:2120448],tree_1[1412627:1409616],tree_1[1415639:1412628]);
csa_3012 csau_3012_i235(A[2126471:2123460],A[2129483:2126472],A[2132495:2129484],tree_1[1418651:1415640],tree_1[1421663:1418652]);
csa_3012 csau_3012_i236(A[2135507:2132496],A[2138519:2135508],A[2141531:2138520],tree_1[1424675:1421664],tree_1[1427687:1424676]);
csa_3012 csau_3012_i237(A[2144543:2141532],A[2147555:2144544],A[2150567:2147556],tree_1[1430699:1427688],tree_1[1433711:1430700]);
csa_3012 csau_3012_i238(A[2153579:2150568],A[2156591:2153580],A[2159603:2156592],tree_1[1436723:1433712],tree_1[1439735:1436724]);
csa_3012 csau_3012_i239(A[2162615:2159604],A[2165627:2162616],A[2168639:2165628],tree_1[1442747:1439736],tree_1[1445759:1442748]);
csa_3012 csau_3012_i240(A[2171651:2168640],A[2174663:2171652],A[2177675:2174664],tree_1[1448771:1445760],tree_1[1451783:1448772]);
csa_3012 csau_3012_i241(A[2180687:2177676],A[2183699:2180688],A[2186711:2183700],tree_1[1454795:1451784],tree_1[1457807:1454796]);
csa_3012 csau_3012_i242(A[2189723:2186712],A[2192735:2189724],A[2195747:2192736],tree_1[1460819:1457808],tree_1[1463831:1460820]);
csa_3012 csau_3012_i243(A[2198759:2195748],A[2201771:2198760],A[2204783:2201772],tree_1[1466843:1463832],tree_1[1469855:1466844]);
csa_3012 csau_3012_i244(A[2207795:2204784],A[2210807:2207796],A[2213819:2210808],tree_1[1472867:1469856],tree_1[1475879:1472868]);
csa_3012 csau_3012_i245(A[2216831:2213820],A[2219843:2216832],A[2222855:2219844],tree_1[1478891:1475880],tree_1[1481903:1478892]);
csa_3012 csau_3012_i246(A[2225867:2222856],A[2228879:2225868],A[2231891:2228880],tree_1[1484915:1481904],tree_1[1487927:1484916]);
csa_3012 csau_3012_i247(A[2234903:2231892],A[2237915:2234904],A[2240927:2237916],tree_1[1490939:1487928],tree_1[1493951:1490940]);
csa_3012 csau_3012_i248(A[2243939:2240928],A[2246951:2243940],A[2249963:2246952],tree_1[1496963:1493952],tree_1[1499975:1496964]);
csa_3012 csau_3012_i249(A[2252975:2249964],A[2255987:2252976],A[2258999:2255988],tree_1[1502987:1499976],tree_1[1505999:1502988]);
csa_3012 csau_3012_i250(A[2262011:2259000],A[2265023:2262012],A[2268035:2265024],tree_1[1509011:1506000],tree_1[1512023:1509012]);
csa_3012 csau_3012_i251(A[2271047:2268036],A[2274059:2271048],A[2277071:2274060],tree_1[1515035:1512024],tree_1[1518047:1515036]);
csa_3012 csau_3012_i252(A[2280083:2277072],A[2283095:2280084],A[2286107:2283096],tree_1[1521059:1518048],tree_1[1524071:1521060]);
csa_3012 csau_3012_i253(A[2289119:2286108],A[2292131:2289120],A[2295143:2292132],tree_1[1527083:1524072],tree_1[1530095:1527084]);
csa_3012 csau_3012_i254(A[2298155:2295144],A[2301167:2298156],A[2304179:2301168],tree_1[1533107:1530096],tree_1[1536119:1533108]);
csa_3012 csau_3012_i255(A[2307191:2304180],A[2310203:2307192],A[2313215:2310204],tree_1[1539131:1536120],tree_1[1542143:1539132]);
csa_3012 csau_3012_i256(A[2316227:2313216],A[2319239:2316228],A[2322251:2319240],tree_1[1545155:1542144],tree_1[1548167:1545156]);
csa_3012 csau_3012_i257(A[2325263:2322252],A[2328275:2325264],A[2331287:2328276],tree_1[1551179:1548168],tree_1[1554191:1551180]);
csa_3012 csau_3012_i258(A[2334299:2331288],A[2337311:2334300],A[2340323:2337312],tree_1[1557203:1554192],tree_1[1560215:1557204]);
csa_3012 csau_3012_i259(A[2343335:2340324],A[2346347:2343336],A[2349359:2346348],tree_1[1563227:1560216],tree_1[1566239:1563228]);
csa_3012 csau_3012_i260(A[2352371:2349360],A[2355383:2352372],A[2358395:2355384],tree_1[1569251:1566240],tree_1[1572263:1569252]);
csa_3012 csau_3012_i261(A[2361407:2358396],A[2364419:2361408],A[2367431:2364420],tree_1[1575275:1572264],tree_1[1578287:1575276]);
csa_3012 csau_3012_i262(A[2370443:2367432],A[2373455:2370444],A[2376467:2373456],tree_1[1581299:1578288],tree_1[1584311:1581300]);
csa_3012 csau_3012_i263(A[2379479:2376468],A[2382491:2379480],A[2385503:2382492],tree_1[1587323:1584312],tree_1[1590335:1587324]);
csa_3012 csau_3012_i264(A[2388515:2385504],A[2391527:2388516],A[2394539:2391528],tree_1[1593347:1590336],tree_1[1596359:1593348]);
csa_3012 csau_3012_i265(A[2397551:2394540],A[2400563:2397552],A[2403575:2400564],tree_1[1599371:1596360],tree_1[1602383:1599372]);
csa_3012 csau_3012_i266(A[2406587:2403576],A[2409599:2406588],A[2412611:2409600],tree_1[1605395:1602384],tree_1[1608407:1605396]);
csa_3012 csau_3012_i267(A[2415623:2412612],A[2418635:2415624],A[2421647:2418636],tree_1[1611419:1608408],tree_1[1614431:1611420]);
csa_3012 csau_3012_i268(A[2424659:2421648],A[2427671:2424660],A[2430683:2427672],tree_1[1617443:1614432],tree_1[1620455:1617444]);
csa_3012 csau_3012_i269(A[2433695:2430684],A[2436707:2433696],A[2439719:2436708],tree_1[1623467:1620456],tree_1[1626479:1623468]);
csa_3012 csau_3012_i270(A[2442731:2439720],A[2445743:2442732],A[2448755:2445744],tree_1[1629491:1626480],tree_1[1632503:1629492]);
csa_3012 csau_3012_i271(A[2451767:2448756],A[2454779:2451768],A[2457791:2454780],tree_1[1635515:1632504],tree_1[1638527:1635516]);
csa_3012 csau_3012_i272(A[2460803:2457792],A[2463815:2460804],A[2466827:2463816],tree_1[1641539:1638528],tree_1[1644551:1641540]);
csa_3012 csau_3012_i273(A[2469839:2466828],A[2472851:2469840],A[2475863:2472852],tree_1[1647563:1644552],tree_1[1650575:1647564]);
csa_3012 csau_3012_i274(A[2478875:2475864],A[2481887:2478876],A[2484899:2481888],tree_1[1653587:1650576],tree_1[1656599:1653588]);
csa_3012 csau_3012_i275(A[2487911:2484900],A[2490923:2487912],A[2493935:2490924],tree_1[1659611:1656600],tree_1[1662623:1659612]);
csa_3012 csau_3012_i276(A[2496947:2493936],A[2499959:2496948],A[2502971:2499960],tree_1[1665635:1662624],tree_1[1668647:1665636]);
csa_3012 csau_3012_i277(A[2505983:2502972],A[2508995:2505984],A[2512007:2508996],tree_1[1671659:1668648],tree_1[1674671:1671660]);
csa_3012 csau_3012_i278(A[2515019:2512008],A[2518031:2515020],A[2521043:2518032],tree_1[1677683:1674672],tree_1[1680695:1677684]);
csa_3012 csau_3012_i279(A[2524055:2521044],A[2527067:2524056],A[2530079:2527068],tree_1[1683707:1680696],tree_1[1686719:1683708]);
csa_3012 csau_3012_i280(A[2533091:2530080],A[2536103:2533092],A[2539115:2536104],tree_1[1689731:1686720],tree_1[1692743:1689732]);
csa_3012 csau_3012_i281(A[2542127:2539116],A[2545139:2542128],A[2548151:2545140],tree_1[1695755:1692744],tree_1[1698767:1695756]);
csa_3012 csau_3012_i282(A[2551163:2548152],A[2554175:2551164],A[2557187:2554176],tree_1[1701779:1698768],tree_1[1704791:1701780]);
csa_3012 csau_3012_i283(A[2560199:2557188],A[2563211:2560200],A[2566223:2563212],tree_1[1707803:1704792],tree_1[1710815:1707804]);
csa_3012 csau_3012_i284(A[2569235:2566224],A[2572247:2569236],A[2575259:2572248],tree_1[1713827:1710816],tree_1[1716839:1713828]);
csa_3012 csau_3012_i285(A[2578271:2575260],A[2581283:2578272],A[2584295:2581284],tree_1[1719851:1716840],tree_1[1722863:1719852]);
csa_3012 csau_3012_i286(A[2587307:2584296],A[2590319:2587308],A[2593331:2590320],tree_1[1725875:1722864],tree_1[1728887:1725876]);
csa_3012 csau_3012_i287(A[2596343:2593332],A[2599355:2596344],A[2602367:2599356],tree_1[1731899:1728888],tree_1[1734911:1731900]);
csa_3012 csau_3012_i288(A[2605379:2602368],A[2608391:2605380],A[2611403:2608392],tree_1[1737923:1734912],tree_1[1740935:1737924]);
csa_3012 csau_3012_i289(A[2614415:2611404],A[2617427:2614416],A[2620439:2617428],tree_1[1743947:1740936],tree_1[1746959:1743948]);
csa_3012 csau_3012_i290(A[2623451:2620440],A[2626463:2623452],A[2629475:2626464],tree_1[1749971:1746960],tree_1[1752983:1749972]);
csa_3012 csau_3012_i291(A[2632487:2629476],A[2635499:2632488],A[2638511:2635500],tree_1[1755995:1752984],tree_1[1759007:1755996]);
csa_3012 csau_3012_i292(A[2641523:2638512],A[2644535:2641524],A[2647547:2644536],tree_1[1762019:1759008],tree_1[1765031:1762020]);
csa_3012 csau_3012_i293(A[2650559:2647548],A[2653571:2650560],A[2656583:2653572],tree_1[1768043:1765032],tree_1[1771055:1768044]);
csa_3012 csau_3012_i294(A[2659595:2656584],A[2662607:2659596],A[2665619:2662608],tree_1[1774067:1771056],tree_1[1777079:1774068]);
csa_3012 csau_3012_i295(A[2668631:2665620],A[2671643:2668632],A[2674655:2671644],tree_1[1780091:1777080],tree_1[1783103:1780092]);
csa_3012 csau_3012_i296(A[2677667:2674656],A[2680679:2677668],A[2683691:2680680],tree_1[1786115:1783104],tree_1[1789127:1786116]);
csa_3012 csau_3012_i297(A[2686703:2683692],A[2689715:2686704],A[2692727:2689716],tree_1[1792139:1789128],tree_1[1795151:1792140]);
csa_3012 csau_3012_i298(A[2695739:2692728],A[2698751:2695740],A[2701763:2698752],tree_1[1798163:1795152],tree_1[1801175:1798164]);
csa_3012 csau_3012_i299(A[2704775:2701764],A[2707787:2704776],A[2710799:2707788],tree_1[1804187:1801176],tree_1[1807199:1804188]);
csa_3012 csau_3012_i300(A[2713811:2710800],A[2716823:2713812],A[2719835:2716824],tree_1[1810211:1807200],tree_1[1813223:1810212]);
csa_3012 csau_3012_i301(A[2722847:2719836],A[2725859:2722848],A[2728871:2725860],tree_1[1816235:1813224],tree_1[1819247:1816236]);
csa_3012 csau_3012_i302(A[2731883:2728872],A[2734895:2731884],A[2737907:2734896],tree_1[1822259:1819248],tree_1[1825271:1822260]);
csa_3012 csau_3012_i303(A[2740919:2737908],A[2743931:2740920],A[2746943:2743932],tree_1[1828283:1825272],tree_1[1831295:1828284]);
csa_3012 csau_3012_i304(A[2749955:2746944],A[2752967:2749956],A[2755979:2752968],tree_1[1834307:1831296],tree_1[1837319:1834308]);
csa_3012 csau_3012_i305(A[2758991:2755980],A[2762003:2758992],A[2765015:2762004],tree_1[1840331:1837320],tree_1[1843343:1840332]);
csa_3012 csau_3012_i306(A[2768027:2765016],A[2771039:2768028],A[2774051:2771040],tree_1[1846355:1843344],tree_1[1849367:1846356]);
csa_3012 csau_3012_i307(A[2777063:2774052],A[2780075:2777064],A[2783087:2780076],tree_1[1852379:1849368],tree_1[1855391:1852380]);
csa_3012 csau_3012_i308(A[2786099:2783088],A[2789111:2786100],A[2792123:2789112],tree_1[1858403:1855392],tree_1[1861415:1858404]);
csa_3012 csau_3012_i309(A[2795135:2792124],A[2798147:2795136],A[2801159:2798148],tree_1[1864427:1861416],tree_1[1867439:1864428]);
csa_3012 csau_3012_i310(A[2804171:2801160],A[2807183:2804172],A[2810195:2807184],tree_1[1870451:1867440],tree_1[1873463:1870452]);
csa_3012 csau_3012_i311(A[2813207:2810196],A[2816219:2813208],A[2819231:2816220],tree_1[1876475:1873464],tree_1[1879487:1876476]);
csa_3012 csau_3012_i312(A[2822243:2819232],A[2825255:2822244],A[2828267:2825256],tree_1[1882499:1879488],tree_1[1885511:1882500]);
csa_3012 csau_3012_i313(A[2831279:2828268],A[2834291:2831280],A[2837303:2834292],tree_1[1888523:1885512],tree_1[1891535:1888524]);
csa_3012 csau_3012_i314(A[2840315:2837304],A[2843327:2840316],A[2846339:2843328],tree_1[1894547:1891536],tree_1[1897559:1894548]);
csa_3012 csau_3012_i315(A[2849351:2846340],A[2852363:2849352],A[2855375:2852364],tree_1[1900571:1897560],tree_1[1903583:1900572]);
csa_3012 csau_3012_i316(A[2858387:2855376],A[2861399:2858388],A[2864411:2861400],tree_1[1906595:1903584],tree_1[1909607:1906596]);
csa_3012 csau_3012_i317(A[2867423:2864412],A[2870435:2867424],A[2873447:2870436],tree_1[1912619:1909608],tree_1[1915631:1912620]);
csa_3012 csau_3012_i318(A[2876459:2873448],A[2879471:2876460],A[2882483:2879472],tree_1[1918643:1915632],tree_1[1921655:1918644]);
csa_3012 csau_3012_i319(A[2885495:2882484],A[2888507:2885496],A[2891519:2888508],tree_1[1924667:1921656],tree_1[1927679:1924668]);
csa_3012 csau_3012_i320(A[2894531:2891520],A[2897543:2894532],A[2900555:2897544],tree_1[1930691:1927680],tree_1[1933703:1930692]);
csa_3012 csau_3012_i321(A[2903567:2900556],A[2906579:2903568],A[2909591:2906580],tree_1[1936715:1933704],tree_1[1939727:1936716]);
csa_3012 csau_3012_i322(A[2912603:2909592],A[2915615:2912604],A[2918627:2915616],tree_1[1942739:1939728],tree_1[1945751:1942740]);
csa_3012 csau_3012_i323(A[2921639:2918628],A[2924651:2921640],A[2927663:2924652],tree_1[1948763:1945752],tree_1[1951775:1948764]);
csa_3012 csau_3012_i324(A[2930675:2927664],A[2933687:2930676],A[2936699:2933688],tree_1[1954787:1951776],tree_1[1957799:1954788]);
csa_3012 csau_3012_i325(A[2939711:2936700],A[2942723:2939712],A[2945735:2942724],tree_1[1960811:1957800],tree_1[1963823:1960812]);
csa_3012 csau_3012_i326(A[2948747:2945736],A[2951759:2948748],A[2954771:2951760],tree_1[1966835:1963824],tree_1[1969847:1966836]);
csa_3012 csau_3012_i327(A[2957783:2954772],A[2960795:2957784],A[2963807:2960796],tree_1[1972859:1969848],tree_1[1975871:1972860]);
csa_3012 csau_3012_i328(A[2966819:2963808],A[2969831:2966820],A[2972843:2969832],tree_1[1978883:1975872],tree_1[1981895:1978884]);
csa_3012 csau_3012_i329(A[2975855:2972844],A[2978867:2975856],A[2981879:2978868],tree_1[1984907:1981896],tree_1[1987919:1984908]);
csa_3012 csau_3012_i330(A[2984891:2981880],A[2987903:2984892],A[2990915:2987904],tree_1[1990931:1987920],tree_1[1993943:1990932]);
csa_3012 csau_3012_i331(A[2993927:2990916],A[2996939:2993928],A[2999951:2996940],tree_1[1996955:1993944],tree_1[1999967:1996956]);
csa_3012 csau_3012_i332(A[3002963:2999952],A[3005975:3002964],A[3008987:3005976],tree_1[2002979:1999968],tree_1[2005991:2002980]);
csa_3012 csau_3012_i333(A[3011999:3008988],A[3015011:3012000],A[3018023:3015012],tree_1[2009003:2005992],tree_1[2012015:2009004]);
csa_3012 csau_3012_i334(A[3021035:3018024],A[3024047:3021036],A[3027059:3024048],tree_1[2015027:2012016],tree_1[2018039:2015028]);
csa_3012 csau_3012_i335(A[3030071:3027060],A[3033083:3030072],A[3036095:3033084],tree_1[2021051:2018040],tree_1[2024063:2021052]);
csa_3012 csau_3012_i336(A[3039107:3036096],A[3042119:3039108],A[3045131:3042120],tree_1[2027075:2024064],tree_1[2030087:2027076]);
csa_3012 csau_3012_i337(A[3048143:3045132],A[3051155:3048144],A[3054167:3051156],tree_1[2033099:2030088],tree_1[2036111:2033100]);
csa_3012 csau_3012_i338(A[3057179:3054168],A[3060191:3057180],A[3063203:3060192],tree_1[2039123:2036112],tree_1[2042135:2039124]);
csa_3012 csau_3012_i339(A[3066215:3063204],A[3069227:3066216],A[3072239:3069228],tree_1[2045147:2042136],tree_1[2048159:2045148]);
csa_3012 csau_3012_i340(A[3075251:3072240],A[3078263:3075252],A[3081275:3078264],tree_1[2051171:2048160],tree_1[2054183:2051172]);
csa_3012 csau_3012_i341(A[3084287:3081276],A[3087299:3084288],A[3090311:3087300],tree_1[2057195:2054184],tree_1[2060207:2057196]);
csa_3012 csau_3012_i342(A[3093323:3090312],A[3096335:3093324],A[3099347:3096336],tree_1[2063219:2060208],tree_1[2066231:2063220]);
csa_3012 csau_3012_i343(A[3102359:3099348],A[3105371:3102360],A[3108383:3105372],tree_1[2069243:2066232],tree_1[2072255:2069244]);
csa_3012 csau_3012_i344(A[3111395:3108384],A[3114407:3111396],A[3117419:3114408],tree_1[2075267:2072256],tree_1[2078279:2075268]);
csa_3012 csau_3012_i345(A[3120431:3117420],A[3123443:3120432],A[3126455:3123444],tree_1[2081291:2078280],tree_1[2084303:2081292]);
csa_3012 csau_3012_i346(A[3129467:3126456],A[3132479:3129468],A[3135491:3132480],tree_1[2087315:2084304],tree_1[2090327:2087316]);
csa_3012 csau_3012_i347(A[3138503:3135492],A[3141515:3138504],A[3144527:3141516],tree_1[2093339:2090328],tree_1[2096351:2093340]);
csa_3012 csau_3012_i348(A[3147539:3144528],A[3150551:3147540],A[3153563:3150552],tree_1[2099363:2096352],tree_1[2102375:2099364]);
csa_3012 csau_3012_i349(A[3156575:3153564],A[3159587:3156576],A[3162599:3159588],tree_1[2105387:2102376],tree_1[2108399:2105388]);
csa_3012 csau_3012_i350(A[3165611:3162600],A[3168623:3165612],A[3171635:3168624],tree_1[2111411:2108400],tree_1[2114423:2111412]);
csa_3012 csau_3012_i351(A[3174647:3171636],A[3177659:3174648],A[3180671:3177660],tree_1[2117435:2114424],tree_1[2120447:2117436]);
csa_3012 csau_3012_i352(A[3183683:3180672],A[3186695:3183684],A[3189707:3186696],tree_1[2123459:2120448],tree_1[2126471:2123460]);
csa_3012 csau_3012_i353(A[3192719:3189708],A[3195731:3192720],A[3198743:3195732],tree_1[2129483:2126472],tree_1[2132495:2129484]);
csa_3012 csau_3012_i354(A[3201755:3198744],A[3204767:3201756],A[3207779:3204768],tree_1[2135507:2132496],tree_1[2138519:2135508]);
csa_3012 csau_3012_i355(A[3210791:3207780],A[3213803:3210792],A[3216815:3213804],tree_1[2141531:2138520],tree_1[2144543:2141532]);
csa_3012 csau_3012_i356(A[3219827:3216816],A[3222839:3219828],A[3225851:3222840],tree_1[2147555:2144544],tree_1[2150567:2147556]);
csa_3012 csau_3012_i357(A[3228863:3225852],A[3231875:3228864],A[3234887:3231876],tree_1[2153579:2150568],tree_1[2156591:2153580]);
csa_3012 csau_3012_i358(A[3237899:3234888],A[3240911:3237900],A[3243923:3240912],tree_1[2159603:2156592],tree_1[2162615:2159604]);
csa_3012 csau_3012_i359(A[3246935:3243924],A[3249947:3246936],A[3252959:3249948],tree_1[2165627:2162616],tree_1[2168639:2165628]);
csa_3012 csau_3012_i360(A[3255971:3252960],A[3258983:3255972],A[3261995:3258984],tree_1[2171651:2168640],tree_1[2174663:2171652]);
csa_3012 csau_3012_i361(A[3265007:3261996],A[3268019:3265008],A[3271031:3268020],tree_1[2177675:2174664],tree_1[2180687:2177676]);
csa_3012 csau_3012_i362(A[3274043:3271032],A[3277055:3274044],A[3280067:3277056],tree_1[2183699:2180688],tree_1[2186711:2183700]);
csa_3012 csau_3012_i363(A[3283079:3280068],A[3286091:3283080],A[3289103:3286092],tree_1[2189723:2186712],tree_1[2192735:2189724]);
csa_3012 csau_3012_i364(A[3292115:3289104],A[3295127:3292116],A[3298139:3295128],tree_1[2195747:2192736],tree_1[2198759:2195748]);
csa_3012 csau_3012_i365(A[3301151:3298140],A[3304163:3301152],A[3307175:3304164],tree_1[2201771:2198760],tree_1[2204783:2201772]);
csa_3012 csau_3012_i366(A[3310187:3307176],A[3313199:3310188],A[3316211:3313200],tree_1[2207795:2204784],tree_1[2210807:2207796]);
csa_3012 csau_3012_i367(A[3319223:3316212],A[3322235:3319224],A[3325247:3322236],tree_1[2213819:2210808],tree_1[2216831:2213820]);
csa_3012 csau_3012_i368(A[3328259:3325248],A[3331271:3328260],A[3334283:3331272],tree_1[2219843:2216832],tree_1[2222855:2219844]);
csa_3012 csau_3012_i369(A[3337295:3334284],A[3340307:3337296],A[3343319:3340308],tree_1[2225867:2222856],tree_1[2228879:2225868]);
csa_3012 csau_3012_i370(A[3346331:3343320],A[3349343:3346332],A[3352355:3349344],tree_1[2231891:2228880],tree_1[2234903:2231892]);
csa_3012 csau_3012_i371(A[3355367:3352356],A[3358379:3355368],A[3361391:3358380],tree_1[2237915:2234904],tree_1[2240927:2237916]);
csa_3012 csau_3012_i372(A[3364403:3361392],A[3367415:3364404],A[3370427:3367416],tree_1[2243939:2240928],tree_1[2246951:2243940]);
csa_3012 csau_3012_i373(A[3373439:3370428],A[3376451:3373440],A[3379463:3376452],tree_1[2249963:2246952],tree_1[2252975:2249964]);
csa_3012 csau_3012_i374(A[3382475:3379464],A[3385487:3382476],A[3388499:3385488],tree_1[2255987:2252976],tree_1[2258999:2255988]);
csa_3012 csau_3012_i375(A[3391511:3388500],A[3394523:3391512],A[3397535:3394524],tree_1[2262011:2259000],tree_1[2265023:2262012]);
csa_3012 csau_3012_i376(A[3400547:3397536],A[3403559:3400548],A[3406571:3403560],tree_1[2268035:2265024],tree_1[2271047:2268036]);
csa_3012 csau_3012_i377(A[3409583:3406572],A[3412595:3409584],A[3415607:3412596],tree_1[2274059:2271048],tree_1[2277071:2274060]);
csa_3012 csau_3012_i378(A[3418619:3415608],A[3421631:3418620],A[3424643:3421632],tree_1[2280083:2277072],tree_1[2283095:2280084]);
csa_3012 csau_3012_i379(A[3427655:3424644],A[3430667:3427656],A[3433679:3430668],tree_1[2286107:2283096],tree_1[2289119:2286108]);
csa_3012 csau_3012_i380(A[3436691:3433680],A[3439703:3436692],A[3442715:3439704],tree_1[2292131:2289120],tree_1[2295143:2292132]);
csa_3012 csau_3012_i381(A[3445727:3442716],A[3448739:3445728],A[3451751:3448740],tree_1[2298155:2295144],tree_1[2301167:2298156]);
csa_3012 csau_3012_i382(A[3454763:3451752],A[3457775:3454764],A[3460787:3457776],tree_1[2304179:2301168],tree_1[2307191:2304180]);
csa_3012 csau_3012_i383(A[3463799:3460788],A[3466811:3463800],A[3469823:3466812],tree_1[2310203:2307192],tree_1[2313215:2310204]);
csa_3012 csau_3012_i384(A[3472835:3469824],A[3475847:3472836],A[3478859:3475848],tree_1[2316227:2313216],tree_1[2319239:2316228]);
csa_3012 csau_3012_i385(A[3481871:3478860],A[3484883:3481872],A[3487895:3484884],tree_1[2322251:2319240],tree_1[2325263:2322252]);
csa_3012 csau_3012_i386(A[3490907:3487896],A[3493919:3490908],A[3496931:3493920],tree_1[2328275:2325264],tree_1[2331287:2328276]);
csa_3012 csau_3012_i387(A[3499943:3496932],A[3502955:3499944],A[3505967:3502956],tree_1[2334299:2331288],tree_1[2337311:2334300]);
csa_3012 csau_3012_i388(A[3508979:3505968],A[3511991:3508980],A[3515003:3511992],tree_1[2340323:2337312],tree_1[2343335:2340324]);
csa_3012 csau_3012_i389(A[3518015:3515004],A[3521027:3518016],A[3524039:3521028],tree_1[2346347:2343336],tree_1[2349359:2346348]);
csa_3012 csau_3012_i390(A[3527051:3524040],A[3530063:3527052],A[3533075:3530064],tree_1[2352371:2349360],tree_1[2355383:2352372]);
csa_3012 csau_3012_i391(A[3536087:3533076],A[3539099:3536088],A[3542111:3539100],tree_1[2358395:2355384],tree_1[2361407:2358396]);
csa_3012 csau_3012_i392(A[3545123:3542112],A[3548135:3545124],A[3551147:3548136],tree_1[2364419:2361408],tree_1[2367431:2364420]);
csa_3012 csau_3012_i393(A[3554159:3551148],A[3557171:3554160],A[3560183:3557172],tree_1[2370443:2367432],tree_1[2373455:2370444]);
csa_3012 csau_3012_i394(A[3563195:3560184],A[3566207:3563196],A[3569219:3566208],tree_1[2376467:2373456],tree_1[2379479:2376468]);
csa_3012 csau_3012_i395(A[3572231:3569220],A[3575243:3572232],A[3578255:3575244],tree_1[2382491:2379480],tree_1[2385503:2382492]);
csa_3012 csau_3012_i396(A[3581267:3578256],A[3584279:3581268],A[3587291:3584280],tree_1[2388515:2385504],tree_1[2391527:2388516]);
csa_3012 csau_3012_i397(A[3590303:3587292],A[3593315:3590304],A[3596327:3593316],tree_1[2394539:2391528],tree_1[2397551:2394540]);
csa_3012 csau_3012_i398(A[3599339:3596328],A[3602351:3599340],A[3605363:3602352],tree_1[2400563:2397552],tree_1[2403575:2400564]);
csa_3012 csau_3012_i399(A[3608375:3605364],A[3611387:3608376],A[3614399:3611388],tree_1[2406587:2403576],tree_1[2409599:2406588]);
csa_3012 csau_3012_i400(A[3617411:3614400],A[3620423:3617412],A[3623435:3620424],tree_1[2412611:2409600],tree_1[2415623:2412612]);
csa_3012 csau_3012_i401(A[3626447:3623436],A[3629459:3626448],A[3632471:3629460],tree_1[2418635:2415624],tree_1[2421647:2418636]);
csa_3012 csau_3012_i402(A[3635483:3632472],A[3638495:3635484],A[3641507:3638496],tree_1[2424659:2421648],tree_1[2427671:2424660]);
csa_3012 csau_3012_i403(A[3644519:3641508],A[3647531:3644520],A[3650543:3647532],tree_1[2430683:2427672],tree_1[2433695:2430684]);
csa_3012 csau_3012_i404(A[3653555:3650544],A[3656567:3653556],A[3659579:3656568],tree_1[2436707:2433696],tree_1[2439719:2436708]);
csa_3012 csau_3012_i405(A[3662591:3659580],A[3665603:3662592],A[3668615:3665604],tree_1[2442731:2439720],tree_1[2445743:2442732]);
csa_3012 csau_3012_i406(A[3671627:3668616],A[3674639:3671628],A[3677651:3674640],tree_1[2448755:2445744],tree_1[2451767:2448756]);
csa_3012 csau_3012_i407(A[3680663:3677652],A[3683675:3680664],A[3686687:3683676],tree_1[2454779:2451768],tree_1[2457791:2454780]);
csa_3012 csau_3012_i408(A[3689699:3686688],A[3692711:3689700],A[3695723:3692712],tree_1[2460803:2457792],tree_1[2463815:2460804]);
csa_3012 csau_3012_i409(A[3698735:3695724],A[3701747:3698736],A[3704759:3701748],tree_1[2466827:2463816],tree_1[2469839:2466828]);
csa_3012 csau_3012_i410(A[3707771:3704760],A[3710783:3707772],A[3713795:3710784],tree_1[2472851:2469840],tree_1[2475863:2472852]);
csa_3012 csau_3012_i411(A[3716807:3713796],A[3719819:3716808],A[3722831:3719820],tree_1[2478875:2475864],tree_1[2481887:2478876]);
csa_3012 csau_3012_i412(A[3725843:3722832],A[3728855:3725844],A[3731867:3728856],tree_1[2484899:2481888],tree_1[2487911:2484900]);
csa_3012 csau_3012_i413(A[3734879:3731868],A[3737891:3734880],A[3740903:3737892],tree_1[2490923:2487912],tree_1[2493935:2490924]);
csa_3012 csau_3012_i414(A[3743915:3740904],A[3746927:3743916],A[3749939:3746928],tree_1[2496947:2493936],tree_1[2499959:2496948]);
csa_3012 csau_3012_i415(A[3752951:3749940],A[3755963:3752952],A[3758975:3755964],tree_1[2502971:2499960],tree_1[2505983:2502972]);
csa_3012 csau_3012_i416(A[3761987:3758976],A[3764999:3761988],A[3768011:3765000],tree_1[2508995:2505984],tree_1[2512007:2508996]);
csa_3012 csau_3012_i417(A[3771023:3768012],A[3774035:3771024],A[3777047:3774036],tree_1[2515019:2512008],tree_1[2518031:2515020]);
csa_3012 csau_3012_i418(A[3780059:3777048],A[3783071:3780060],A[3786083:3783072],tree_1[2521043:2518032],tree_1[2524055:2521044]);
csa_3012 csau_3012_i419(A[3789095:3786084],A[3792107:3789096],A[3795119:3792108],tree_1[2527067:2524056],tree_1[2530079:2527068]);
csa_3012 csau_3012_i420(A[3798131:3795120],A[3801143:3798132],A[3804155:3801144],tree_1[2533091:2530080],tree_1[2536103:2533092]);
csa_3012 csau_3012_i421(A[3807167:3804156],A[3810179:3807168],A[3813191:3810180],tree_1[2539115:2536104],tree_1[2542127:2539116]);
csa_3012 csau_3012_i422(A[3816203:3813192],A[3819215:3816204],A[3822227:3819216],tree_1[2545139:2542128],tree_1[2548151:2545140]);
csa_3012 csau_3012_i423(A[3825239:3822228],A[3828251:3825240],A[3831263:3828252],tree_1[2551163:2548152],tree_1[2554175:2551164]);
csa_3012 csau_3012_i424(A[3834275:3831264],A[3837287:3834276],A[3840299:3837288],tree_1[2557187:2554176],tree_1[2560199:2557188]);
csa_3012 csau_3012_i425(A[3843311:3840300],A[3846323:3843312],A[3849335:3846324],tree_1[2563211:2560200],tree_1[2566223:2563212]);
csa_3012 csau_3012_i426(A[3852347:3849336],A[3855359:3852348],A[3858371:3855360],tree_1[2569235:2566224],tree_1[2572247:2569236]);
csa_3012 csau_3012_i427(A[3861383:3858372],A[3864395:3861384],A[3867407:3864396],tree_1[2575259:2572248],tree_1[2578271:2575260]);
csa_3012 csau_3012_i428(A[3870419:3867408],A[3873431:3870420],A[3876443:3873432],tree_1[2581283:2578272],tree_1[2584295:2581284]);
csa_3012 csau_3012_i429(A[3879455:3876444],A[3882467:3879456],A[3885479:3882468],tree_1[2587307:2584296],tree_1[2590319:2587308]);
csa_3012 csau_3012_i430(A[3888491:3885480],A[3891503:3888492],A[3894515:3891504],tree_1[2593331:2590320],tree_1[2596343:2593332]);
csa_3012 csau_3012_i431(A[3897527:3894516],A[3900539:3897528],A[3903551:3900540],tree_1[2599355:2596344],tree_1[2602367:2599356]);
csa_3012 csau_3012_i432(A[3906563:3903552],A[3909575:3906564],A[3912587:3909576],tree_1[2605379:2602368],tree_1[2608391:2605380]);
csa_3012 csau_3012_i433(A[3915599:3912588],A[3918611:3915600],A[3921623:3918612],tree_1[2611403:2608392],tree_1[2614415:2611404]);
csa_3012 csau_3012_i434(A[3924635:3921624],A[3927647:3924636],A[3930659:3927648],tree_1[2617427:2614416],tree_1[2620439:2617428]);
csa_3012 csau_3012_i435(A[3933671:3930660],A[3936683:3933672],A[3939695:3936684],tree_1[2623451:2620440],tree_1[2626463:2623452]);
csa_3012 csau_3012_i436(A[3942707:3939696],A[3945719:3942708],A[3948731:3945720],tree_1[2629475:2626464],tree_1[2632487:2629476]);
csa_3012 csau_3012_i437(A[3951743:3948732],A[3954755:3951744],A[3957767:3954756],tree_1[2635499:2632488],tree_1[2638511:2635500]);
csa_3012 csau_3012_i438(A[3960779:3957768],A[3963791:3960780],A[3966803:3963792],tree_1[2641523:2638512],tree_1[2644535:2641524]);
csa_3012 csau_3012_i439(A[3969815:3966804],A[3972827:3969816],A[3975839:3972828],tree_1[2647547:2644536],tree_1[2650559:2647548]);
csa_3012 csau_3012_i440(A[3978851:3975840],A[3981863:3978852],A[3984875:3981864],tree_1[2653571:2650560],tree_1[2656583:2653572]);
csa_3012 csau_3012_i441(A[3987887:3984876],A[3990899:3987888],A[3993911:3990900],tree_1[2659595:2656584],tree_1[2662607:2659596]);
csa_3012 csau_3012_i442(A[3996923:3993912],A[3999935:3996924],A[4002947:3999936],tree_1[2665619:2662608],tree_1[2668631:2665620]);
csa_3012 csau_3012_i443(A[4005959:4002948],A[4008971:4005960],A[4011983:4008972],tree_1[2671643:2668632],tree_1[2674655:2671644]);
csa_3012 csau_3012_i444(A[4014995:4011984],A[4018007:4014996],A[4021019:4018008],tree_1[2677667:2674656],tree_1[2680679:2677668]);
csa_3012 csau_3012_i445(A[4024031:4021020],A[4027043:4024032],A[4030055:4027044],tree_1[2683691:2680680],tree_1[2686703:2683692]);
csa_3012 csau_3012_i446(A[4033067:4030056],A[4036079:4033068],A[4039091:4036080],tree_1[2689715:2686704],tree_1[2692727:2689716]);
csa_3012 csau_3012_i447(A[4042103:4039092],A[4045115:4042104],A[4048127:4045116],tree_1[2695739:2692728],tree_1[2698751:2695740]);
csa_3012 csau_3012_i448(A[4051139:4048128],A[4054151:4051140],A[4057163:4054152],tree_1[2701763:2698752],tree_1[2704775:2701764]);
csa_3012 csau_3012_i449(A[4060175:4057164],A[4063187:4060176],A[4066199:4063188],tree_1[2707787:2704776],tree_1[2710799:2707788]);
csa_3012 csau_3012_i450(A[4069211:4066200],A[4072223:4069212],A[4075235:4072224],tree_1[2713811:2710800],tree_1[2716823:2713812]);
csa_3012 csau_3012_i451(A[4078247:4075236],A[4081259:4078248],A[4084271:4081260],tree_1[2719835:2716824],tree_1[2722847:2719836]);
csa_3012 csau_3012_i452(A[4087283:4084272],A[4090295:4087284],A[4093307:4090296],tree_1[2725859:2722848],tree_1[2728871:2725860]);
csa_3012 csau_3012_i453(A[4096319:4093308],A[4099331:4096320],A[4102343:4099332],tree_1[2731883:2728872],tree_1[2734895:2731884]);
csa_3012 csau_3012_i454(A[4105355:4102344],A[4108367:4105356],A[4111379:4108368],tree_1[2737907:2734896],tree_1[2740919:2737908]);
csa_3012 csau_3012_i455(A[4114391:4111380],A[4117403:4114392],A[4120415:4117404],tree_1[2743931:2740920],tree_1[2746943:2743932]);
csa_3012 csau_3012_i456(A[4123427:4120416],A[4126439:4123428],A[4129451:4126440],tree_1[2749955:2746944],tree_1[2752967:2749956]);
csa_3012 csau_3012_i457(A[4132463:4129452],A[4135475:4132464],A[4138487:4135476],tree_1[2755979:2752968],tree_1[2758991:2755980]);
csa_3012 csau_3012_i458(A[4141499:4138488],A[4144511:4141500],A[4147523:4144512],tree_1[2762003:2758992],tree_1[2765015:2762004]);
csa_3012 csau_3012_i459(A[4150535:4147524],A[4153547:4150536],A[4156559:4153548],tree_1[2768027:2765016],tree_1[2771039:2768028]);
csa_3012 csau_3012_i460(A[4159571:4156560],A[4162583:4159572],A[4165595:4162584],tree_1[2774051:2771040],tree_1[2777063:2774052]);
csa_3012 csau_3012_i461(A[4168607:4165596],A[4171619:4168608],A[4174631:4171620],tree_1[2780075:2777064],tree_1[2783087:2780076]);
csa_3012 csau_3012_i462(A[4177643:4174632],A[4180655:4177644],A[4183667:4180656],tree_1[2786099:2783088],tree_1[2789111:2786100]);
csa_3012 csau_3012_i463(A[4186679:4183668],A[4189691:4186680],A[4192703:4189692],tree_1[2792123:2789112],tree_1[2795135:2792124]);
csa_3012 csau_3012_i464(A[4195715:4192704],A[4198727:4195716],A[4201739:4198728],tree_1[2798147:2795136],tree_1[2801159:2798148]);
csa_3012 csau_3012_i465(A[4204751:4201740],A[4207763:4204752],A[4210775:4207764],tree_1[2804171:2801160],tree_1[2807183:2804172]);
csa_3012 csau_3012_i466(A[4213787:4210776],A[4216799:4213788],A[4219811:4216800],tree_1[2810195:2807184],tree_1[2813207:2810196]);
csa_3012 csau_3012_i467(A[4222823:4219812],A[4225835:4222824],A[4228847:4225836],tree_1[2816219:2813208],tree_1[2819231:2816220]);
csa_3012 csau_3012_i468(A[4231859:4228848],A[4234871:4231860],A[4237883:4234872],tree_1[2822243:2819232],tree_1[2825255:2822244]);
csa_3012 csau_3012_i469(A[4240895:4237884],A[4243907:4240896],A[4246919:4243908],tree_1[2828267:2825256],tree_1[2831279:2828268]);
csa_3012 csau_3012_i470(A[4249931:4246920],A[4252943:4249932],A[4255955:4252944],tree_1[2834291:2831280],tree_1[2837303:2834292]);
csa_3012 csau_3012_i471(A[4258967:4255956],A[4261979:4258968],A[4264991:4261980],tree_1[2840315:2837304],tree_1[2843327:2840316]);
csa_3012 csau_3012_i472(A[4268003:4264992],A[4271015:4268004],A[4274027:4271016],tree_1[2846339:2843328],tree_1[2849351:2846340]);
csa_3012 csau_3012_i473(A[4277039:4274028],A[4280051:4277040],A[4283063:4280052],tree_1[2852363:2849352],tree_1[2855375:2852364]);
csa_3012 csau_3012_i474(A[4286075:4283064],A[4289087:4286076],A[4292099:4289088],tree_1[2858387:2855376],tree_1[2861399:2858388]);
csa_3012 csau_3012_i475(A[4295111:4292100],A[4298123:4295112],A[4301135:4298124],tree_1[2864411:2861400],tree_1[2867423:2864412]);
csa_3012 csau_3012_i476(A[4304147:4301136],A[4307159:4304148],A[4310171:4307160],tree_1[2870435:2867424],tree_1[2873447:2870436]);
csa_3012 csau_3012_i477(A[4313183:4310172],A[4316195:4313184],A[4319207:4316196],tree_1[2876459:2873448],tree_1[2879471:2876460]);
csa_3012 csau_3012_i478(A[4322219:4319208],A[4325231:4322220],A[4328243:4325232],tree_1[2882483:2879472],tree_1[2885495:2882484]);
csa_3012 csau_3012_i479(A[4331255:4328244],A[4334267:4331256],A[4337279:4334268],tree_1[2888507:2885496],tree_1[2891519:2888508]);
csa_3012 csau_3012_i480(A[4340291:4337280],A[4343303:4340292],A[4346315:4343304],tree_1[2894531:2891520],tree_1[2897543:2894532]);
csa_3012 csau_3012_i481(A[4349327:4346316],A[4352339:4349328],A[4355351:4352340],tree_1[2900555:2897544],tree_1[2903567:2900556]);
csa_3012 csau_3012_i482(A[4358363:4355352],A[4361375:4358364],A[4364387:4361376],tree_1[2906579:2903568],tree_1[2909591:2906580]);
csa_3012 csau_3012_i483(A[4367399:4364388],A[4370411:4367400],A[4373423:4370412],tree_1[2912603:2909592],tree_1[2915615:2912604]);
csa_3012 csau_3012_i484(A[4376435:4373424],A[4379447:4376436],A[4382459:4379448],tree_1[2918627:2915616],tree_1[2921639:2918628]);
csa_3012 csau_3012_i485(A[4385471:4382460],A[4388483:4385472],A[4391495:4388484],tree_1[2924651:2921640],tree_1[2927663:2924652]);
csa_3012 csau_3012_i486(A[4394507:4391496],A[4397519:4394508],A[4400531:4397520],tree_1[2930675:2927664],tree_1[2933687:2930676]);
csa_3012 csau_3012_i487(A[4403543:4400532],A[4406555:4403544],A[4409567:4406556],tree_1[2936699:2933688],tree_1[2939711:2936700]);
csa_3012 csau_3012_i488(A[4412579:4409568],A[4415591:4412580],A[4418603:4415592],tree_1[2942723:2939712],tree_1[2945735:2942724]);
csa_3012 csau_3012_i489(A[4421615:4418604],A[4424627:4421616],A[4427639:4424628],tree_1[2948747:2945736],tree_1[2951759:2948748]);
csa_3012 csau_3012_i490(A[4430651:4427640],A[4433663:4430652],A[4436675:4433664],tree_1[2954771:2951760],tree_1[2957783:2954772]);
csa_3012 csau_3012_i491(A[4439687:4436676],A[4442699:4439688],A[4445711:4442700],tree_1[2960795:2957784],tree_1[2963807:2960796]);
csa_3012 csau_3012_i492(A[4448723:4445712],A[4451735:4448724],A[4454747:4451736],tree_1[2966819:2963808],tree_1[2969831:2966820]);
csa_3012 csau_3012_i493(A[4457759:4454748],A[4460771:4457760],A[4463783:4460772],tree_1[2972843:2969832],tree_1[2975855:2972844]);
csa_3012 csau_3012_i494(A[4466795:4463784],A[4469807:4466796],A[4472819:4469808],tree_1[2978867:2975856],tree_1[2981879:2978868]);
csa_3012 csau_3012_i495(A[4475831:4472820],A[4478843:4475832],A[4481855:4478844],tree_1[2984891:2981880],tree_1[2987903:2984892]);
csa_3012 csau_3012_i496(A[4484867:4481856],A[4487879:4484868],A[4490891:4487880],tree_1[2990915:2987904],tree_1[2993927:2990916]);
csa_3012 csau_3012_i497(A[4493903:4490892],A[4496915:4493904],A[4499927:4496916],tree_1[2996939:2993928],tree_1[2999951:2996940]);
csa_3012 csau_3012_i498(A[4502939:4499928],A[4505951:4502940],A[4508963:4505952],tree_1[3002963:2999952],tree_1[3005975:3002964]);
csa_3012 csau_3012_i499(A[4511975:4508964],A[4514987:4511976],A[4517999:4514988],tree_1[3008987:3005976],tree_1[3011999:3008988]);
csa_3012 csau_3012_i500(A[4521011:4518000],A[4524023:4521012],A[4527035:4524024],tree_1[3015011:3012000],tree_1[3018023:3015012]);
csa_3012 csau_3012_i501(A[4530047:4527036],A[4533059:4530048],A[4536071:4533060],tree_1[3021035:3018024],tree_1[3024047:3021036]);
// layer-2
csa_3012 csau_3012_i502(tree_1[3011:0],tree_1[6023:3012],tree_1[9035:6024],tree_2[3011:0],tree_2[6023:3012]);
csa_3012 csau_3012_i503(tree_1[12047:9036],tree_1[15059:12048],tree_1[18071:15060],tree_2[9035:6024],tree_2[12047:9036]);
csa_3012 csau_3012_i504(tree_1[21083:18072],tree_1[24095:21084],tree_1[27107:24096],tree_2[15059:12048],tree_2[18071:15060]);
csa_3012 csau_3012_i505(tree_1[30119:27108],tree_1[33131:30120],tree_1[36143:33132],tree_2[21083:18072],tree_2[24095:21084]);
csa_3012 csau_3012_i506(tree_1[39155:36144],tree_1[42167:39156],tree_1[45179:42168],tree_2[27107:24096],tree_2[30119:27108]);
csa_3012 csau_3012_i507(tree_1[48191:45180],tree_1[51203:48192],tree_1[54215:51204],tree_2[33131:30120],tree_2[36143:33132]);
csa_3012 csau_3012_i508(tree_1[57227:54216],tree_1[60239:57228],tree_1[63251:60240],tree_2[39155:36144],tree_2[42167:39156]);
csa_3012 csau_3012_i509(tree_1[66263:63252],tree_1[69275:66264],tree_1[72287:69276],tree_2[45179:42168],tree_2[48191:45180]);
csa_3012 csau_3012_i510(tree_1[75299:72288],tree_1[78311:75300],tree_1[81323:78312],tree_2[51203:48192],tree_2[54215:51204]);
csa_3012 csau_3012_i511(tree_1[84335:81324],tree_1[87347:84336],tree_1[90359:87348],tree_2[57227:54216],tree_2[60239:57228]);
csa_3012 csau_3012_i512(tree_1[93371:90360],tree_1[96383:93372],tree_1[99395:96384],tree_2[63251:60240],tree_2[66263:63252]);
csa_3012 csau_3012_i513(tree_1[102407:99396],tree_1[105419:102408],tree_1[108431:105420],tree_2[69275:66264],tree_2[72287:69276]);
csa_3012 csau_3012_i514(tree_1[111443:108432],tree_1[114455:111444],tree_1[117467:114456],tree_2[75299:72288],tree_2[78311:75300]);
csa_3012 csau_3012_i515(tree_1[120479:117468],tree_1[123491:120480],tree_1[126503:123492],tree_2[81323:78312],tree_2[84335:81324]);
csa_3012 csau_3012_i516(tree_1[129515:126504],tree_1[132527:129516],tree_1[135539:132528],tree_2[87347:84336],tree_2[90359:87348]);
csa_3012 csau_3012_i517(tree_1[138551:135540],tree_1[141563:138552],tree_1[144575:141564],tree_2[93371:90360],tree_2[96383:93372]);
csa_3012 csau_3012_i518(tree_1[147587:144576],tree_1[150599:147588],tree_1[153611:150600],tree_2[99395:96384],tree_2[102407:99396]);
csa_3012 csau_3012_i519(tree_1[156623:153612],tree_1[159635:156624],tree_1[162647:159636],tree_2[105419:102408],tree_2[108431:105420]);
csa_3012 csau_3012_i520(tree_1[165659:162648],tree_1[168671:165660],tree_1[171683:168672],tree_2[111443:108432],tree_2[114455:111444]);
csa_3012 csau_3012_i521(tree_1[174695:171684],tree_1[177707:174696],tree_1[180719:177708],tree_2[117467:114456],tree_2[120479:117468]);
csa_3012 csau_3012_i522(tree_1[183731:180720],tree_1[186743:183732],tree_1[189755:186744],tree_2[123491:120480],tree_2[126503:123492]);
csa_3012 csau_3012_i523(tree_1[192767:189756],tree_1[195779:192768],tree_1[198791:195780],tree_2[129515:126504],tree_2[132527:129516]);
csa_3012 csau_3012_i524(tree_1[201803:198792],tree_1[204815:201804],tree_1[207827:204816],tree_2[135539:132528],tree_2[138551:135540]);
csa_3012 csau_3012_i525(tree_1[210839:207828],tree_1[213851:210840],tree_1[216863:213852],tree_2[141563:138552],tree_2[144575:141564]);
csa_3012 csau_3012_i526(tree_1[219875:216864],tree_1[222887:219876],tree_1[225899:222888],tree_2[147587:144576],tree_2[150599:147588]);
csa_3012 csau_3012_i527(tree_1[228911:225900],tree_1[231923:228912],tree_1[234935:231924],tree_2[153611:150600],tree_2[156623:153612]);
csa_3012 csau_3012_i528(tree_1[237947:234936],tree_1[240959:237948],tree_1[243971:240960],tree_2[159635:156624],tree_2[162647:159636]);
csa_3012 csau_3012_i529(tree_1[246983:243972],tree_1[249995:246984],tree_1[253007:249996],tree_2[165659:162648],tree_2[168671:165660]);
csa_3012 csau_3012_i530(tree_1[256019:253008],tree_1[259031:256020],tree_1[262043:259032],tree_2[171683:168672],tree_2[174695:171684]);
csa_3012 csau_3012_i531(tree_1[265055:262044],tree_1[268067:265056],tree_1[271079:268068],tree_2[177707:174696],tree_2[180719:177708]);
csa_3012 csau_3012_i532(tree_1[274091:271080],tree_1[277103:274092],tree_1[280115:277104],tree_2[183731:180720],tree_2[186743:183732]);
csa_3012 csau_3012_i533(tree_1[283127:280116],tree_1[286139:283128],tree_1[289151:286140],tree_2[189755:186744],tree_2[192767:189756]);
csa_3012 csau_3012_i534(tree_1[292163:289152],tree_1[295175:292164],tree_1[298187:295176],tree_2[195779:192768],tree_2[198791:195780]);
csa_3012 csau_3012_i535(tree_1[301199:298188],tree_1[304211:301200],tree_1[307223:304212],tree_2[201803:198792],tree_2[204815:201804]);
csa_3012 csau_3012_i536(tree_1[310235:307224],tree_1[313247:310236],tree_1[316259:313248],tree_2[207827:204816],tree_2[210839:207828]);
csa_3012 csau_3012_i537(tree_1[319271:316260],tree_1[322283:319272],tree_1[325295:322284],tree_2[213851:210840],tree_2[216863:213852]);
csa_3012 csau_3012_i538(tree_1[328307:325296],tree_1[331319:328308],tree_1[334331:331320],tree_2[219875:216864],tree_2[222887:219876]);
csa_3012 csau_3012_i539(tree_1[337343:334332],tree_1[340355:337344],tree_1[343367:340356],tree_2[225899:222888],tree_2[228911:225900]);
csa_3012 csau_3012_i540(tree_1[346379:343368],tree_1[349391:346380],tree_1[352403:349392],tree_2[231923:228912],tree_2[234935:231924]);
csa_3012 csau_3012_i541(tree_1[355415:352404],tree_1[358427:355416],tree_1[361439:358428],tree_2[237947:234936],tree_2[240959:237948]);
csa_3012 csau_3012_i542(tree_1[364451:361440],tree_1[367463:364452],tree_1[370475:367464],tree_2[243971:240960],tree_2[246983:243972]);
csa_3012 csau_3012_i543(tree_1[373487:370476],tree_1[376499:373488],tree_1[379511:376500],tree_2[249995:246984],tree_2[253007:249996]);
csa_3012 csau_3012_i544(tree_1[382523:379512],tree_1[385535:382524],tree_1[388547:385536],tree_2[256019:253008],tree_2[259031:256020]);
csa_3012 csau_3012_i545(tree_1[391559:388548],tree_1[394571:391560],tree_1[397583:394572],tree_2[262043:259032],tree_2[265055:262044]);
csa_3012 csau_3012_i546(tree_1[400595:397584],tree_1[403607:400596],tree_1[406619:403608],tree_2[268067:265056],tree_2[271079:268068]);
csa_3012 csau_3012_i547(tree_1[409631:406620],tree_1[412643:409632],tree_1[415655:412644],tree_2[274091:271080],tree_2[277103:274092]);
csa_3012 csau_3012_i548(tree_1[418667:415656],tree_1[421679:418668],tree_1[424691:421680],tree_2[280115:277104],tree_2[283127:280116]);
csa_3012 csau_3012_i549(tree_1[427703:424692],tree_1[430715:427704],tree_1[433727:430716],tree_2[286139:283128],tree_2[289151:286140]);
csa_3012 csau_3012_i550(tree_1[436739:433728],tree_1[439751:436740],tree_1[442763:439752],tree_2[292163:289152],tree_2[295175:292164]);
csa_3012 csau_3012_i551(tree_1[445775:442764],tree_1[448787:445776],tree_1[451799:448788],tree_2[298187:295176],tree_2[301199:298188]);
csa_3012 csau_3012_i552(tree_1[454811:451800],tree_1[457823:454812],tree_1[460835:457824],tree_2[304211:301200],tree_2[307223:304212]);
csa_3012 csau_3012_i553(tree_1[463847:460836],tree_1[466859:463848],tree_1[469871:466860],tree_2[310235:307224],tree_2[313247:310236]);
csa_3012 csau_3012_i554(tree_1[472883:469872],tree_1[475895:472884],tree_1[478907:475896],tree_2[316259:313248],tree_2[319271:316260]);
csa_3012 csau_3012_i555(tree_1[481919:478908],tree_1[484931:481920],tree_1[487943:484932],tree_2[322283:319272],tree_2[325295:322284]);
csa_3012 csau_3012_i556(tree_1[490955:487944],tree_1[493967:490956],tree_1[496979:493968],tree_2[328307:325296],tree_2[331319:328308]);
csa_3012 csau_3012_i557(tree_1[499991:496980],tree_1[503003:499992],tree_1[506015:503004],tree_2[334331:331320],tree_2[337343:334332]);
csa_3012 csau_3012_i558(tree_1[509027:506016],tree_1[512039:509028],tree_1[515051:512040],tree_2[340355:337344],tree_2[343367:340356]);
csa_3012 csau_3012_i559(tree_1[518063:515052],tree_1[521075:518064],tree_1[524087:521076],tree_2[346379:343368],tree_2[349391:346380]);
csa_3012 csau_3012_i560(tree_1[527099:524088],tree_1[530111:527100],tree_1[533123:530112],tree_2[352403:349392],tree_2[355415:352404]);
csa_3012 csau_3012_i561(tree_1[536135:533124],tree_1[539147:536136],tree_1[542159:539148],tree_2[358427:355416],tree_2[361439:358428]);
csa_3012 csau_3012_i562(tree_1[545171:542160],tree_1[548183:545172],tree_1[551195:548184],tree_2[364451:361440],tree_2[367463:364452]);
csa_3012 csau_3012_i563(tree_1[554207:551196],tree_1[557219:554208],tree_1[560231:557220],tree_2[370475:367464],tree_2[373487:370476]);
csa_3012 csau_3012_i564(tree_1[563243:560232],tree_1[566255:563244],tree_1[569267:566256],tree_2[376499:373488],tree_2[379511:376500]);
csa_3012 csau_3012_i565(tree_1[572279:569268],tree_1[575291:572280],tree_1[578303:575292],tree_2[382523:379512],tree_2[385535:382524]);
csa_3012 csau_3012_i566(tree_1[581315:578304],tree_1[584327:581316],tree_1[587339:584328],tree_2[388547:385536],tree_2[391559:388548]);
csa_3012 csau_3012_i567(tree_1[590351:587340],tree_1[593363:590352],tree_1[596375:593364],tree_2[394571:391560],tree_2[397583:394572]);
csa_3012 csau_3012_i568(tree_1[599387:596376],tree_1[602399:599388],tree_1[605411:602400],tree_2[400595:397584],tree_2[403607:400596]);
csa_3012 csau_3012_i569(tree_1[608423:605412],tree_1[611435:608424],tree_1[614447:611436],tree_2[406619:403608],tree_2[409631:406620]);
csa_3012 csau_3012_i570(tree_1[617459:614448],tree_1[620471:617460],tree_1[623483:620472],tree_2[412643:409632],tree_2[415655:412644]);
csa_3012 csau_3012_i571(tree_1[626495:623484],tree_1[629507:626496],tree_1[632519:629508],tree_2[418667:415656],tree_2[421679:418668]);
csa_3012 csau_3012_i572(tree_1[635531:632520],tree_1[638543:635532],tree_1[641555:638544],tree_2[424691:421680],tree_2[427703:424692]);
csa_3012 csau_3012_i573(tree_1[644567:641556],tree_1[647579:644568],tree_1[650591:647580],tree_2[430715:427704],tree_2[433727:430716]);
csa_3012 csau_3012_i574(tree_1[653603:650592],tree_1[656615:653604],tree_1[659627:656616],tree_2[436739:433728],tree_2[439751:436740]);
csa_3012 csau_3012_i575(tree_1[662639:659628],tree_1[665651:662640],tree_1[668663:665652],tree_2[442763:439752],tree_2[445775:442764]);
csa_3012 csau_3012_i576(tree_1[671675:668664],tree_1[674687:671676],tree_1[677699:674688],tree_2[448787:445776],tree_2[451799:448788]);
csa_3012 csau_3012_i577(tree_1[680711:677700],tree_1[683723:680712],tree_1[686735:683724],tree_2[454811:451800],tree_2[457823:454812]);
csa_3012 csau_3012_i578(tree_1[689747:686736],tree_1[692759:689748],tree_1[695771:692760],tree_2[460835:457824],tree_2[463847:460836]);
csa_3012 csau_3012_i579(tree_1[698783:695772],tree_1[701795:698784],tree_1[704807:701796],tree_2[466859:463848],tree_2[469871:466860]);
csa_3012 csau_3012_i580(tree_1[707819:704808],tree_1[710831:707820],tree_1[713843:710832],tree_2[472883:469872],tree_2[475895:472884]);
csa_3012 csau_3012_i581(tree_1[716855:713844],tree_1[719867:716856],tree_1[722879:719868],tree_2[478907:475896],tree_2[481919:478908]);
csa_3012 csau_3012_i582(tree_1[725891:722880],tree_1[728903:725892],tree_1[731915:728904],tree_2[484931:481920],tree_2[487943:484932]);
csa_3012 csau_3012_i583(tree_1[734927:731916],tree_1[737939:734928],tree_1[740951:737940],tree_2[490955:487944],tree_2[493967:490956]);
csa_3012 csau_3012_i584(tree_1[743963:740952],tree_1[746975:743964],tree_1[749987:746976],tree_2[496979:493968],tree_2[499991:496980]);
csa_3012 csau_3012_i585(tree_1[752999:749988],tree_1[756011:753000],tree_1[759023:756012],tree_2[503003:499992],tree_2[506015:503004]);
csa_3012 csau_3012_i586(tree_1[762035:759024],tree_1[765047:762036],tree_1[768059:765048],tree_2[509027:506016],tree_2[512039:509028]);
csa_3012 csau_3012_i587(tree_1[771071:768060],tree_1[774083:771072],tree_1[777095:774084],tree_2[515051:512040],tree_2[518063:515052]);
csa_3012 csau_3012_i588(tree_1[780107:777096],tree_1[783119:780108],tree_1[786131:783120],tree_2[521075:518064],tree_2[524087:521076]);
csa_3012 csau_3012_i589(tree_1[789143:786132],tree_1[792155:789144],tree_1[795167:792156],tree_2[527099:524088],tree_2[530111:527100]);
csa_3012 csau_3012_i590(tree_1[798179:795168],tree_1[801191:798180],tree_1[804203:801192],tree_2[533123:530112],tree_2[536135:533124]);
csa_3012 csau_3012_i591(tree_1[807215:804204],tree_1[810227:807216],tree_1[813239:810228],tree_2[539147:536136],tree_2[542159:539148]);
csa_3012 csau_3012_i592(tree_1[816251:813240],tree_1[819263:816252],tree_1[822275:819264],tree_2[545171:542160],tree_2[548183:545172]);
csa_3012 csau_3012_i593(tree_1[825287:822276],tree_1[828299:825288],tree_1[831311:828300],tree_2[551195:548184],tree_2[554207:551196]);
csa_3012 csau_3012_i594(tree_1[834323:831312],tree_1[837335:834324],tree_1[840347:837336],tree_2[557219:554208],tree_2[560231:557220]);
csa_3012 csau_3012_i595(tree_1[843359:840348],tree_1[846371:843360],tree_1[849383:846372],tree_2[563243:560232],tree_2[566255:563244]);
csa_3012 csau_3012_i596(tree_1[852395:849384],tree_1[855407:852396],tree_1[858419:855408],tree_2[569267:566256],tree_2[572279:569268]);
csa_3012 csau_3012_i597(tree_1[861431:858420],tree_1[864443:861432],tree_1[867455:864444],tree_2[575291:572280],tree_2[578303:575292]);
csa_3012 csau_3012_i598(tree_1[870467:867456],tree_1[873479:870468],tree_1[876491:873480],tree_2[581315:578304],tree_2[584327:581316]);
csa_3012 csau_3012_i599(tree_1[879503:876492],tree_1[882515:879504],tree_1[885527:882516],tree_2[587339:584328],tree_2[590351:587340]);
csa_3012 csau_3012_i600(tree_1[888539:885528],tree_1[891551:888540],tree_1[894563:891552],tree_2[593363:590352],tree_2[596375:593364]);
csa_3012 csau_3012_i601(tree_1[897575:894564],tree_1[900587:897576],tree_1[903599:900588],tree_2[599387:596376],tree_2[602399:599388]);
csa_3012 csau_3012_i602(tree_1[906611:903600],tree_1[909623:906612],tree_1[912635:909624],tree_2[605411:602400],tree_2[608423:605412]);
csa_3012 csau_3012_i603(tree_1[915647:912636],tree_1[918659:915648],tree_1[921671:918660],tree_2[611435:608424],tree_2[614447:611436]);
csa_3012 csau_3012_i604(tree_1[924683:921672],tree_1[927695:924684],tree_1[930707:927696],tree_2[617459:614448],tree_2[620471:617460]);
csa_3012 csau_3012_i605(tree_1[933719:930708],tree_1[936731:933720],tree_1[939743:936732],tree_2[623483:620472],tree_2[626495:623484]);
csa_3012 csau_3012_i606(tree_1[942755:939744],tree_1[945767:942756],tree_1[948779:945768],tree_2[629507:626496],tree_2[632519:629508]);
csa_3012 csau_3012_i607(tree_1[951791:948780],tree_1[954803:951792],tree_1[957815:954804],tree_2[635531:632520],tree_2[638543:635532]);
csa_3012 csau_3012_i608(tree_1[960827:957816],tree_1[963839:960828],tree_1[966851:963840],tree_2[641555:638544],tree_2[644567:641556]);
csa_3012 csau_3012_i609(tree_1[969863:966852],tree_1[972875:969864],tree_1[975887:972876],tree_2[647579:644568],tree_2[650591:647580]);
csa_3012 csau_3012_i610(tree_1[978899:975888],tree_1[981911:978900],tree_1[984923:981912],tree_2[653603:650592],tree_2[656615:653604]);
csa_3012 csau_3012_i611(tree_1[987935:984924],tree_1[990947:987936],tree_1[993959:990948],tree_2[659627:656616],tree_2[662639:659628]);
csa_3012 csau_3012_i612(tree_1[996971:993960],tree_1[999983:996972],tree_1[1002995:999984],tree_2[665651:662640],tree_2[668663:665652]);
csa_3012 csau_3012_i613(tree_1[1006007:1002996],tree_1[1009019:1006008],tree_1[1012031:1009020],tree_2[671675:668664],tree_2[674687:671676]);
csa_3012 csau_3012_i614(tree_1[1015043:1012032],tree_1[1018055:1015044],tree_1[1021067:1018056],tree_2[677699:674688],tree_2[680711:677700]);
csa_3012 csau_3012_i615(tree_1[1024079:1021068],tree_1[1027091:1024080],tree_1[1030103:1027092],tree_2[683723:680712],tree_2[686735:683724]);
csa_3012 csau_3012_i616(tree_1[1033115:1030104],tree_1[1036127:1033116],tree_1[1039139:1036128],tree_2[689747:686736],tree_2[692759:689748]);
csa_3012 csau_3012_i617(tree_1[1042151:1039140],tree_1[1045163:1042152],tree_1[1048175:1045164],tree_2[695771:692760],tree_2[698783:695772]);
csa_3012 csau_3012_i618(tree_1[1051187:1048176],tree_1[1054199:1051188],tree_1[1057211:1054200],tree_2[701795:698784],tree_2[704807:701796]);
csa_3012 csau_3012_i619(tree_1[1060223:1057212],tree_1[1063235:1060224],tree_1[1066247:1063236],tree_2[707819:704808],tree_2[710831:707820]);
csa_3012 csau_3012_i620(tree_1[1069259:1066248],tree_1[1072271:1069260],tree_1[1075283:1072272],tree_2[713843:710832],tree_2[716855:713844]);
csa_3012 csau_3012_i621(tree_1[1078295:1075284],tree_1[1081307:1078296],tree_1[1084319:1081308],tree_2[719867:716856],tree_2[722879:719868]);
csa_3012 csau_3012_i622(tree_1[1087331:1084320],tree_1[1090343:1087332],tree_1[1093355:1090344],tree_2[725891:722880],tree_2[728903:725892]);
csa_3012 csau_3012_i623(tree_1[1096367:1093356],tree_1[1099379:1096368],tree_1[1102391:1099380],tree_2[731915:728904],tree_2[734927:731916]);
csa_3012 csau_3012_i624(tree_1[1105403:1102392],tree_1[1108415:1105404],tree_1[1111427:1108416],tree_2[737939:734928],tree_2[740951:737940]);
csa_3012 csau_3012_i625(tree_1[1114439:1111428],tree_1[1117451:1114440],tree_1[1120463:1117452],tree_2[743963:740952],tree_2[746975:743964]);
csa_3012 csau_3012_i626(tree_1[1123475:1120464],tree_1[1126487:1123476],tree_1[1129499:1126488],tree_2[749987:746976],tree_2[752999:749988]);
csa_3012 csau_3012_i627(tree_1[1132511:1129500],tree_1[1135523:1132512],tree_1[1138535:1135524],tree_2[756011:753000],tree_2[759023:756012]);
csa_3012 csau_3012_i628(tree_1[1141547:1138536],tree_1[1144559:1141548],tree_1[1147571:1144560],tree_2[762035:759024],tree_2[765047:762036]);
csa_3012 csau_3012_i629(tree_1[1150583:1147572],tree_1[1153595:1150584],tree_1[1156607:1153596],tree_2[768059:765048],tree_2[771071:768060]);
csa_3012 csau_3012_i630(tree_1[1159619:1156608],tree_1[1162631:1159620],tree_1[1165643:1162632],tree_2[774083:771072],tree_2[777095:774084]);
csa_3012 csau_3012_i631(tree_1[1168655:1165644],tree_1[1171667:1168656],tree_1[1174679:1171668],tree_2[780107:777096],tree_2[783119:780108]);
csa_3012 csau_3012_i632(tree_1[1177691:1174680],tree_1[1180703:1177692],tree_1[1183715:1180704],tree_2[786131:783120],tree_2[789143:786132]);
csa_3012 csau_3012_i633(tree_1[1186727:1183716],tree_1[1189739:1186728],tree_1[1192751:1189740],tree_2[792155:789144],tree_2[795167:792156]);
csa_3012 csau_3012_i634(tree_1[1195763:1192752],tree_1[1198775:1195764],tree_1[1201787:1198776],tree_2[798179:795168],tree_2[801191:798180]);
csa_3012 csau_3012_i635(tree_1[1204799:1201788],tree_1[1207811:1204800],tree_1[1210823:1207812],tree_2[804203:801192],tree_2[807215:804204]);
csa_3012 csau_3012_i636(tree_1[1213835:1210824],tree_1[1216847:1213836],tree_1[1219859:1216848],tree_2[810227:807216],tree_2[813239:810228]);
csa_3012 csau_3012_i637(tree_1[1222871:1219860],tree_1[1225883:1222872],tree_1[1228895:1225884],tree_2[816251:813240],tree_2[819263:816252]);
csa_3012 csau_3012_i638(tree_1[1231907:1228896],tree_1[1234919:1231908],tree_1[1237931:1234920],tree_2[822275:819264],tree_2[825287:822276]);
csa_3012 csau_3012_i639(tree_1[1240943:1237932],tree_1[1243955:1240944],tree_1[1246967:1243956],tree_2[828299:825288],tree_2[831311:828300]);
csa_3012 csau_3012_i640(tree_1[1249979:1246968],tree_1[1252991:1249980],tree_1[1256003:1252992],tree_2[834323:831312],tree_2[837335:834324]);
csa_3012 csau_3012_i641(tree_1[1259015:1256004],tree_1[1262027:1259016],tree_1[1265039:1262028],tree_2[840347:837336],tree_2[843359:840348]);
csa_3012 csau_3012_i642(tree_1[1268051:1265040],tree_1[1271063:1268052],tree_1[1274075:1271064],tree_2[846371:843360],tree_2[849383:846372]);
csa_3012 csau_3012_i643(tree_1[1277087:1274076],tree_1[1280099:1277088],tree_1[1283111:1280100],tree_2[852395:849384],tree_2[855407:852396]);
csa_3012 csau_3012_i644(tree_1[1286123:1283112],tree_1[1289135:1286124],tree_1[1292147:1289136],tree_2[858419:855408],tree_2[861431:858420]);
csa_3012 csau_3012_i645(tree_1[1295159:1292148],tree_1[1298171:1295160],tree_1[1301183:1298172],tree_2[864443:861432],tree_2[867455:864444]);
csa_3012 csau_3012_i646(tree_1[1304195:1301184],tree_1[1307207:1304196],tree_1[1310219:1307208],tree_2[870467:867456],tree_2[873479:870468]);
csa_3012 csau_3012_i647(tree_1[1313231:1310220],tree_1[1316243:1313232],tree_1[1319255:1316244],tree_2[876491:873480],tree_2[879503:876492]);
csa_3012 csau_3012_i648(tree_1[1322267:1319256],tree_1[1325279:1322268],tree_1[1328291:1325280],tree_2[882515:879504],tree_2[885527:882516]);
csa_3012 csau_3012_i649(tree_1[1331303:1328292],tree_1[1334315:1331304],tree_1[1337327:1334316],tree_2[888539:885528],tree_2[891551:888540]);
csa_3012 csau_3012_i650(tree_1[1340339:1337328],tree_1[1343351:1340340],tree_1[1346363:1343352],tree_2[894563:891552],tree_2[897575:894564]);
csa_3012 csau_3012_i651(tree_1[1349375:1346364],tree_1[1352387:1349376],tree_1[1355399:1352388],tree_2[900587:897576],tree_2[903599:900588]);
csa_3012 csau_3012_i652(tree_1[1358411:1355400],tree_1[1361423:1358412],tree_1[1364435:1361424],tree_2[906611:903600],tree_2[909623:906612]);
csa_3012 csau_3012_i653(tree_1[1367447:1364436],tree_1[1370459:1367448],tree_1[1373471:1370460],tree_2[912635:909624],tree_2[915647:912636]);
csa_3012 csau_3012_i654(tree_1[1376483:1373472],tree_1[1379495:1376484],tree_1[1382507:1379496],tree_2[918659:915648],tree_2[921671:918660]);
csa_3012 csau_3012_i655(tree_1[1385519:1382508],tree_1[1388531:1385520],tree_1[1391543:1388532],tree_2[924683:921672],tree_2[927695:924684]);
csa_3012 csau_3012_i656(tree_1[1394555:1391544],tree_1[1397567:1394556],tree_1[1400579:1397568],tree_2[930707:927696],tree_2[933719:930708]);
csa_3012 csau_3012_i657(tree_1[1403591:1400580],tree_1[1406603:1403592],tree_1[1409615:1406604],tree_2[936731:933720],tree_2[939743:936732]);
csa_3012 csau_3012_i658(tree_1[1412627:1409616],tree_1[1415639:1412628],tree_1[1418651:1415640],tree_2[942755:939744],tree_2[945767:942756]);
csa_3012 csau_3012_i659(tree_1[1421663:1418652],tree_1[1424675:1421664],tree_1[1427687:1424676],tree_2[948779:945768],tree_2[951791:948780]);
csa_3012 csau_3012_i660(tree_1[1430699:1427688],tree_1[1433711:1430700],tree_1[1436723:1433712],tree_2[954803:951792],tree_2[957815:954804]);
csa_3012 csau_3012_i661(tree_1[1439735:1436724],tree_1[1442747:1439736],tree_1[1445759:1442748],tree_2[960827:957816],tree_2[963839:960828]);
csa_3012 csau_3012_i662(tree_1[1448771:1445760],tree_1[1451783:1448772],tree_1[1454795:1451784],tree_2[966851:963840],tree_2[969863:966852]);
csa_3012 csau_3012_i663(tree_1[1457807:1454796],tree_1[1460819:1457808],tree_1[1463831:1460820],tree_2[972875:969864],tree_2[975887:972876]);
csa_3012 csau_3012_i664(tree_1[1466843:1463832],tree_1[1469855:1466844],tree_1[1472867:1469856],tree_2[978899:975888],tree_2[981911:978900]);
csa_3012 csau_3012_i665(tree_1[1475879:1472868],tree_1[1478891:1475880],tree_1[1481903:1478892],tree_2[984923:981912],tree_2[987935:984924]);
csa_3012 csau_3012_i666(tree_1[1484915:1481904],tree_1[1487927:1484916],tree_1[1490939:1487928],tree_2[990947:987936],tree_2[993959:990948]);
csa_3012 csau_3012_i667(tree_1[1493951:1490940],tree_1[1496963:1493952],tree_1[1499975:1496964],tree_2[996971:993960],tree_2[999983:996972]);
csa_3012 csau_3012_i668(tree_1[1502987:1499976],tree_1[1505999:1502988],tree_1[1509011:1506000],tree_2[1002995:999984],tree_2[1006007:1002996]);
csa_3012 csau_3012_i669(tree_1[1512023:1509012],tree_1[1515035:1512024],tree_1[1518047:1515036],tree_2[1009019:1006008],tree_2[1012031:1009020]);
csa_3012 csau_3012_i670(tree_1[1521059:1518048],tree_1[1524071:1521060],tree_1[1527083:1524072],tree_2[1015043:1012032],tree_2[1018055:1015044]);
csa_3012 csau_3012_i671(tree_1[1530095:1527084],tree_1[1533107:1530096],tree_1[1536119:1533108],tree_2[1021067:1018056],tree_2[1024079:1021068]);
csa_3012 csau_3012_i672(tree_1[1539131:1536120],tree_1[1542143:1539132],tree_1[1545155:1542144],tree_2[1027091:1024080],tree_2[1030103:1027092]);
csa_3012 csau_3012_i673(tree_1[1548167:1545156],tree_1[1551179:1548168],tree_1[1554191:1551180],tree_2[1033115:1030104],tree_2[1036127:1033116]);
csa_3012 csau_3012_i674(tree_1[1557203:1554192],tree_1[1560215:1557204],tree_1[1563227:1560216],tree_2[1039139:1036128],tree_2[1042151:1039140]);
csa_3012 csau_3012_i675(tree_1[1566239:1563228],tree_1[1569251:1566240],tree_1[1572263:1569252],tree_2[1045163:1042152],tree_2[1048175:1045164]);
csa_3012 csau_3012_i676(tree_1[1575275:1572264],tree_1[1578287:1575276],tree_1[1581299:1578288],tree_2[1051187:1048176],tree_2[1054199:1051188]);
csa_3012 csau_3012_i677(tree_1[1584311:1581300],tree_1[1587323:1584312],tree_1[1590335:1587324],tree_2[1057211:1054200],tree_2[1060223:1057212]);
csa_3012 csau_3012_i678(tree_1[1593347:1590336],tree_1[1596359:1593348],tree_1[1599371:1596360],tree_2[1063235:1060224],tree_2[1066247:1063236]);
csa_3012 csau_3012_i679(tree_1[1602383:1599372],tree_1[1605395:1602384],tree_1[1608407:1605396],tree_2[1069259:1066248],tree_2[1072271:1069260]);
csa_3012 csau_3012_i680(tree_1[1611419:1608408],tree_1[1614431:1611420],tree_1[1617443:1614432],tree_2[1075283:1072272],tree_2[1078295:1075284]);
csa_3012 csau_3012_i681(tree_1[1620455:1617444],tree_1[1623467:1620456],tree_1[1626479:1623468],tree_2[1081307:1078296],tree_2[1084319:1081308]);
csa_3012 csau_3012_i682(tree_1[1629491:1626480],tree_1[1632503:1629492],tree_1[1635515:1632504],tree_2[1087331:1084320],tree_2[1090343:1087332]);
csa_3012 csau_3012_i683(tree_1[1638527:1635516],tree_1[1641539:1638528],tree_1[1644551:1641540],tree_2[1093355:1090344],tree_2[1096367:1093356]);
csa_3012 csau_3012_i684(tree_1[1647563:1644552],tree_1[1650575:1647564],tree_1[1653587:1650576],tree_2[1099379:1096368],tree_2[1102391:1099380]);
csa_3012 csau_3012_i685(tree_1[1656599:1653588],tree_1[1659611:1656600],tree_1[1662623:1659612],tree_2[1105403:1102392],tree_2[1108415:1105404]);
csa_3012 csau_3012_i686(tree_1[1665635:1662624],tree_1[1668647:1665636],tree_1[1671659:1668648],tree_2[1111427:1108416],tree_2[1114439:1111428]);
csa_3012 csau_3012_i687(tree_1[1674671:1671660],tree_1[1677683:1674672],tree_1[1680695:1677684],tree_2[1117451:1114440],tree_2[1120463:1117452]);
csa_3012 csau_3012_i688(tree_1[1683707:1680696],tree_1[1686719:1683708],tree_1[1689731:1686720],tree_2[1123475:1120464],tree_2[1126487:1123476]);
csa_3012 csau_3012_i689(tree_1[1692743:1689732],tree_1[1695755:1692744],tree_1[1698767:1695756],tree_2[1129499:1126488],tree_2[1132511:1129500]);
csa_3012 csau_3012_i690(tree_1[1701779:1698768],tree_1[1704791:1701780],tree_1[1707803:1704792],tree_2[1135523:1132512],tree_2[1138535:1135524]);
csa_3012 csau_3012_i691(tree_1[1710815:1707804],tree_1[1713827:1710816],tree_1[1716839:1713828],tree_2[1141547:1138536],tree_2[1144559:1141548]);
csa_3012 csau_3012_i692(tree_1[1719851:1716840],tree_1[1722863:1719852],tree_1[1725875:1722864],tree_2[1147571:1144560],tree_2[1150583:1147572]);
csa_3012 csau_3012_i693(tree_1[1728887:1725876],tree_1[1731899:1728888],tree_1[1734911:1731900],tree_2[1153595:1150584],tree_2[1156607:1153596]);
csa_3012 csau_3012_i694(tree_1[1737923:1734912],tree_1[1740935:1737924],tree_1[1743947:1740936],tree_2[1159619:1156608],tree_2[1162631:1159620]);
csa_3012 csau_3012_i695(tree_1[1746959:1743948],tree_1[1749971:1746960],tree_1[1752983:1749972],tree_2[1165643:1162632],tree_2[1168655:1165644]);
csa_3012 csau_3012_i696(tree_1[1755995:1752984],tree_1[1759007:1755996],tree_1[1762019:1759008],tree_2[1171667:1168656],tree_2[1174679:1171668]);
csa_3012 csau_3012_i697(tree_1[1765031:1762020],tree_1[1768043:1765032],tree_1[1771055:1768044],tree_2[1177691:1174680],tree_2[1180703:1177692]);
csa_3012 csau_3012_i698(tree_1[1774067:1771056],tree_1[1777079:1774068],tree_1[1780091:1777080],tree_2[1183715:1180704],tree_2[1186727:1183716]);
csa_3012 csau_3012_i699(tree_1[1783103:1780092],tree_1[1786115:1783104],tree_1[1789127:1786116],tree_2[1189739:1186728],tree_2[1192751:1189740]);
csa_3012 csau_3012_i700(tree_1[1792139:1789128],tree_1[1795151:1792140],tree_1[1798163:1795152],tree_2[1195763:1192752],tree_2[1198775:1195764]);
csa_3012 csau_3012_i701(tree_1[1801175:1798164],tree_1[1804187:1801176],tree_1[1807199:1804188],tree_2[1201787:1198776],tree_2[1204799:1201788]);
csa_3012 csau_3012_i702(tree_1[1810211:1807200],tree_1[1813223:1810212],tree_1[1816235:1813224],tree_2[1207811:1204800],tree_2[1210823:1207812]);
csa_3012 csau_3012_i703(tree_1[1819247:1816236],tree_1[1822259:1819248],tree_1[1825271:1822260],tree_2[1213835:1210824],tree_2[1216847:1213836]);
csa_3012 csau_3012_i704(tree_1[1828283:1825272],tree_1[1831295:1828284],tree_1[1834307:1831296],tree_2[1219859:1216848],tree_2[1222871:1219860]);
csa_3012 csau_3012_i705(tree_1[1837319:1834308],tree_1[1840331:1837320],tree_1[1843343:1840332],tree_2[1225883:1222872],tree_2[1228895:1225884]);
csa_3012 csau_3012_i706(tree_1[1846355:1843344],tree_1[1849367:1846356],tree_1[1852379:1849368],tree_2[1231907:1228896],tree_2[1234919:1231908]);
csa_3012 csau_3012_i707(tree_1[1855391:1852380],tree_1[1858403:1855392],tree_1[1861415:1858404],tree_2[1237931:1234920],tree_2[1240943:1237932]);
csa_3012 csau_3012_i708(tree_1[1864427:1861416],tree_1[1867439:1864428],tree_1[1870451:1867440],tree_2[1243955:1240944],tree_2[1246967:1243956]);
csa_3012 csau_3012_i709(tree_1[1873463:1870452],tree_1[1876475:1873464],tree_1[1879487:1876476],tree_2[1249979:1246968],tree_2[1252991:1249980]);
csa_3012 csau_3012_i710(tree_1[1882499:1879488],tree_1[1885511:1882500],tree_1[1888523:1885512],tree_2[1256003:1252992],tree_2[1259015:1256004]);
csa_3012 csau_3012_i711(tree_1[1891535:1888524],tree_1[1894547:1891536],tree_1[1897559:1894548],tree_2[1262027:1259016],tree_2[1265039:1262028]);
csa_3012 csau_3012_i712(tree_1[1900571:1897560],tree_1[1903583:1900572],tree_1[1906595:1903584],tree_2[1268051:1265040],tree_2[1271063:1268052]);
csa_3012 csau_3012_i713(tree_1[1909607:1906596],tree_1[1912619:1909608],tree_1[1915631:1912620],tree_2[1274075:1271064],tree_2[1277087:1274076]);
csa_3012 csau_3012_i714(tree_1[1918643:1915632],tree_1[1921655:1918644],tree_1[1924667:1921656],tree_2[1280099:1277088],tree_2[1283111:1280100]);
csa_3012 csau_3012_i715(tree_1[1927679:1924668],tree_1[1930691:1927680],tree_1[1933703:1930692],tree_2[1286123:1283112],tree_2[1289135:1286124]);
csa_3012 csau_3012_i716(tree_1[1936715:1933704],tree_1[1939727:1936716],tree_1[1942739:1939728],tree_2[1292147:1289136],tree_2[1295159:1292148]);
csa_3012 csau_3012_i717(tree_1[1945751:1942740],tree_1[1948763:1945752],tree_1[1951775:1948764],tree_2[1298171:1295160],tree_2[1301183:1298172]);
csa_3012 csau_3012_i718(tree_1[1954787:1951776],tree_1[1957799:1954788],tree_1[1960811:1957800],tree_2[1304195:1301184],tree_2[1307207:1304196]);
csa_3012 csau_3012_i719(tree_1[1963823:1960812],tree_1[1966835:1963824],tree_1[1969847:1966836],tree_2[1310219:1307208],tree_2[1313231:1310220]);
csa_3012 csau_3012_i720(tree_1[1972859:1969848],tree_1[1975871:1972860],tree_1[1978883:1975872],tree_2[1316243:1313232],tree_2[1319255:1316244]);
csa_3012 csau_3012_i721(tree_1[1981895:1978884],tree_1[1984907:1981896],tree_1[1987919:1984908],tree_2[1322267:1319256],tree_2[1325279:1322268]);
csa_3012 csau_3012_i722(tree_1[1990931:1987920],tree_1[1993943:1990932],tree_1[1996955:1993944],tree_2[1328291:1325280],tree_2[1331303:1328292]);
csa_3012 csau_3012_i723(tree_1[1999967:1996956],tree_1[2002979:1999968],tree_1[2005991:2002980],tree_2[1334315:1331304],tree_2[1337327:1334316]);
csa_3012 csau_3012_i724(tree_1[2009003:2005992],tree_1[2012015:2009004],tree_1[2015027:2012016],tree_2[1340339:1337328],tree_2[1343351:1340340]);
csa_3012 csau_3012_i725(tree_1[2018039:2015028],tree_1[2021051:2018040],tree_1[2024063:2021052],tree_2[1346363:1343352],tree_2[1349375:1346364]);
csa_3012 csau_3012_i726(tree_1[2027075:2024064],tree_1[2030087:2027076],tree_1[2033099:2030088],tree_2[1352387:1349376],tree_2[1355399:1352388]);
csa_3012 csau_3012_i727(tree_1[2036111:2033100],tree_1[2039123:2036112],tree_1[2042135:2039124],tree_2[1358411:1355400],tree_2[1361423:1358412]);
csa_3012 csau_3012_i728(tree_1[2045147:2042136],tree_1[2048159:2045148],tree_1[2051171:2048160],tree_2[1364435:1361424],tree_2[1367447:1364436]);
csa_3012 csau_3012_i729(tree_1[2054183:2051172],tree_1[2057195:2054184],tree_1[2060207:2057196],tree_2[1370459:1367448],tree_2[1373471:1370460]);
csa_3012 csau_3012_i730(tree_1[2063219:2060208],tree_1[2066231:2063220],tree_1[2069243:2066232],tree_2[1376483:1373472],tree_2[1379495:1376484]);
csa_3012 csau_3012_i731(tree_1[2072255:2069244],tree_1[2075267:2072256],tree_1[2078279:2075268],tree_2[1382507:1379496],tree_2[1385519:1382508]);
csa_3012 csau_3012_i732(tree_1[2081291:2078280],tree_1[2084303:2081292],tree_1[2087315:2084304],tree_2[1388531:1385520],tree_2[1391543:1388532]);
csa_3012 csau_3012_i733(tree_1[2090327:2087316],tree_1[2093339:2090328],tree_1[2096351:2093340],tree_2[1394555:1391544],tree_2[1397567:1394556]);
csa_3012 csau_3012_i734(tree_1[2099363:2096352],tree_1[2102375:2099364],tree_1[2105387:2102376],tree_2[1400579:1397568],tree_2[1403591:1400580]);
csa_3012 csau_3012_i735(tree_1[2108399:2105388],tree_1[2111411:2108400],tree_1[2114423:2111412],tree_2[1406603:1403592],tree_2[1409615:1406604]);
csa_3012 csau_3012_i736(tree_1[2117435:2114424],tree_1[2120447:2117436],tree_1[2123459:2120448],tree_2[1412627:1409616],tree_2[1415639:1412628]);
csa_3012 csau_3012_i737(tree_1[2126471:2123460],tree_1[2129483:2126472],tree_1[2132495:2129484],tree_2[1418651:1415640],tree_2[1421663:1418652]);
csa_3012 csau_3012_i738(tree_1[2135507:2132496],tree_1[2138519:2135508],tree_1[2141531:2138520],tree_2[1424675:1421664],tree_2[1427687:1424676]);
csa_3012 csau_3012_i739(tree_1[2144543:2141532],tree_1[2147555:2144544],tree_1[2150567:2147556],tree_2[1430699:1427688],tree_2[1433711:1430700]);
csa_3012 csau_3012_i740(tree_1[2153579:2150568],tree_1[2156591:2153580],tree_1[2159603:2156592],tree_2[1436723:1433712],tree_2[1439735:1436724]);
csa_3012 csau_3012_i741(tree_1[2162615:2159604],tree_1[2165627:2162616],tree_1[2168639:2165628],tree_2[1442747:1439736],tree_2[1445759:1442748]);
csa_3012 csau_3012_i742(tree_1[2171651:2168640],tree_1[2174663:2171652],tree_1[2177675:2174664],tree_2[1448771:1445760],tree_2[1451783:1448772]);
csa_3012 csau_3012_i743(tree_1[2180687:2177676],tree_1[2183699:2180688],tree_1[2186711:2183700],tree_2[1454795:1451784],tree_2[1457807:1454796]);
csa_3012 csau_3012_i744(tree_1[2189723:2186712],tree_1[2192735:2189724],tree_1[2195747:2192736],tree_2[1460819:1457808],tree_2[1463831:1460820]);
csa_3012 csau_3012_i745(tree_1[2198759:2195748],tree_1[2201771:2198760],tree_1[2204783:2201772],tree_2[1466843:1463832],tree_2[1469855:1466844]);
csa_3012 csau_3012_i746(tree_1[2207795:2204784],tree_1[2210807:2207796],tree_1[2213819:2210808],tree_2[1472867:1469856],tree_2[1475879:1472868]);
csa_3012 csau_3012_i747(tree_1[2216831:2213820],tree_1[2219843:2216832],tree_1[2222855:2219844],tree_2[1478891:1475880],tree_2[1481903:1478892]);
csa_3012 csau_3012_i748(tree_1[2225867:2222856],tree_1[2228879:2225868],tree_1[2231891:2228880],tree_2[1484915:1481904],tree_2[1487927:1484916]);
csa_3012 csau_3012_i749(tree_1[2234903:2231892],tree_1[2237915:2234904],tree_1[2240927:2237916],tree_2[1490939:1487928],tree_2[1493951:1490940]);
csa_3012 csau_3012_i750(tree_1[2243939:2240928],tree_1[2246951:2243940],tree_1[2249963:2246952],tree_2[1496963:1493952],tree_2[1499975:1496964]);
csa_3012 csau_3012_i751(tree_1[2252975:2249964],tree_1[2255987:2252976],tree_1[2258999:2255988],tree_2[1502987:1499976],tree_2[1505999:1502988]);
csa_3012 csau_3012_i752(tree_1[2262011:2259000],tree_1[2265023:2262012],tree_1[2268035:2265024],tree_2[1509011:1506000],tree_2[1512023:1509012]);
csa_3012 csau_3012_i753(tree_1[2271047:2268036],tree_1[2274059:2271048],tree_1[2277071:2274060],tree_2[1515035:1512024],tree_2[1518047:1515036]);
csa_3012 csau_3012_i754(tree_1[2280083:2277072],tree_1[2283095:2280084],tree_1[2286107:2283096],tree_2[1521059:1518048],tree_2[1524071:1521060]);
csa_3012 csau_3012_i755(tree_1[2289119:2286108],tree_1[2292131:2289120],tree_1[2295143:2292132],tree_2[1527083:1524072],tree_2[1530095:1527084]);
csa_3012 csau_3012_i756(tree_1[2298155:2295144],tree_1[2301167:2298156],tree_1[2304179:2301168],tree_2[1533107:1530096],tree_2[1536119:1533108]);
csa_3012 csau_3012_i757(tree_1[2307191:2304180],tree_1[2310203:2307192],tree_1[2313215:2310204],tree_2[1539131:1536120],tree_2[1542143:1539132]);
csa_3012 csau_3012_i758(tree_1[2316227:2313216],tree_1[2319239:2316228],tree_1[2322251:2319240],tree_2[1545155:1542144],tree_2[1548167:1545156]);
csa_3012 csau_3012_i759(tree_1[2325263:2322252],tree_1[2328275:2325264],tree_1[2331287:2328276],tree_2[1551179:1548168],tree_2[1554191:1551180]);
csa_3012 csau_3012_i760(tree_1[2334299:2331288],tree_1[2337311:2334300],tree_1[2340323:2337312],tree_2[1557203:1554192],tree_2[1560215:1557204]);
csa_3012 csau_3012_i761(tree_1[2343335:2340324],tree_1[2346347:2343336],tree_1[2349359:2346348],tree_2[1563227:1560216],tree_2[1566239:1563228]);
csa_3012 csau_3012_i762(tree_1[2352371:2349360],tree_1[2355383:2352372],tree_1[2358395:2355384],tree_2[1569251:1566240],tree_2[1572263:1569252]);
csa_3012 csau_3012_i763(tree_1[2361407:2358396],tree_1[2364419:2361408],tree_1[2367431:2364420],tree_2[1575275:1572264],tree_2[1578287:1575276]);
csa_3012 csau_3012_i764(tree_1[2370443:2367432],tree_1[2373455:2370444],tree_1[2376467:2373456],tree_2[1581299:1578288],tree_2[1584311:1581300]);
csa_3012 csau_3012_i765(tree_1[2379479:2376468],tree_1[2382491:2379480],tree_1[2385503:2382492],tree_2[1587323:1584312],tree_2[1590335:1587324]);
csa_3012 csau_3012_i766(tree_1[2388515:2385504],tree_1[2391527:2388516],tree_1[2394539:2391528],tree_2[1593347:1590336],tree_2[1596359:1593348]);
csa_3012 csau_3012_i767(tree_1[2397551:2394540],tree_1[2400563:2397552],tree_1[2403575:2400564],tree_2[1599371:1596360],tree_2[1602383:1599372]);
csa_3012 csau_3012_i768(tree_1[2406587:2403576],tree_1[2409599:2406588],tree_1[2412611:2409600],tree_2[1605395:1602384],tree_2[1608407:1605396]);
csa_3012 csau_3012_i769(tree_1[2415623:2412612],tree_1[2418635:2415624],tree_1[2421647:2418636],tree_2[1611419:1608408],tree_2[1614431:1611420]);
csa_3012 csau_3012_i770(tree_1[2424659:2421648],tree_1[2427671:2424660],tree_1[2430683:2427672],tree_2[1617443:1614432],tree_2[1620455:1617444]);
csa_3012 csau_3012_i771(tree_1[2433695:2430684],tree_1[2436707:2433696],tree_1[2439719:2436708],tree_2[1623467:1620456],tree_2[1626479:1623468]);
csa_3012 csau_3012_i772(tree_1[2442731:2439720],tree_1[2445743:2442732],tree_1[2448755:2445744],tree_2[1629491:1626480],tree_2[1632503:1629492]);
csa_3012 csau_3012_i773(tree_1[2451767:2448756],tree_1[2454779:2451768],tree_1[2457791:2454780],tree_2[1635515:1632504],tree_2[1638527:1635516]);
csa_3012 csau_3012_i774(tree_1[2460803:2457792],tree_1[2463815:2460804],tree_1[2466827:2463816],tree_2[1641539:1638528],tree_2[1644551:1641540]);
csa_3012 csau_3012_i775(tree_1[2469839:2466828],tree_1[2472851:2469840],tree_1[2475863:2472852],tree_2[1647563:1644552],tree_2[1650575:1647564]);
csa_3012 csau_3012_i776(tree_1[2478875:2475864],tree_1[2481887:2478876],tree_1[2484899:2481888],tree_2[1653587:1650576],tree_2[1656599:1653588]);
csa_3012 csau_3012_i777(tree_1[2487911:2484900],tree_1[2490923:2487912],tree_1[2493935:2490924],tree_2[1659611:1656600],tree_2[1662623:1659612]);
csa_3012 csau_3012_i778(tree_1[2496947:2493936],tree_1[2499959:2496948],tree_1[2502971:2499960],tree_2[1665635:1662624],tree_2[1668647:1665636]);
csa_3012 csau_3012_i779(tree_1[2505983:2502972],tree_1[2508995:2505984],tree_1[2512007:2508996],tree_2[1671659:1668648],tree_2[1674671:1671660]);
csa_3012 csau_3012_i780(tree_1[2515019:2512008],tree_1[2518031:2515020],tree_1[2521043:2518032],tree_2[1677683:1674672],tree_2[1680695:1677684]);
csa_3012 csau_3012_i781(tree_1[2524055:2521044],tree_1[2527067:2524056],tree_1[2530079:2527068],tree_2[1683707:1680696],tree_2[1686719:1683708]);
csa_3012 csau_3012_i782(tree_1[2533091:2530080],tree_1[2536103:2533092],tree_1[2539115:2536104],tree_2[1689731:1686720],tree_2[1692743:1689732]);
csa_3012 csau_3012_i783(tree_1[2542127:2539116],tree_1[2545139:2542128],tree_1[2548151:2545140],tree_2[1695755:1692744],tree_2[1698767:1695756]);
csa_3012 csau_3012_i784(tree_1[2551163:2548152],tree_1[2554175:2551164],tree_1[2557187:2554176],tree_2[1701779:1698768],tree_2[1704791:1701780]);
csa_3012 csau_3012_i785(tree_1[2560199:2557188],tree_1[2563211:2560200],tree_1[2566223:2563212],tree_2[1707803:1704792],tree_2[1710815:1707804]);
csa_3012 csau_3012_i786(tree_1[2569235:2566224],tree_1[2572247:2569236],tree_1[2575259:2572248],tree_2[1713827:1710816],tree_2[1716839:1713828]);
csa_3012 csau_3012_i787(tree_1[2578271:2575260],tree_1[2581283:2578272],tree_1[2584295:2581284],tree_2[1719851:1716840],tree_2[1722863:1719852]);
csa_3012 csau_3012_i788(tree_1[2587307:2584296],tree_1[2590319:2587308],tree_1[2593331:2590320],tree_2[1725875:1722864],tree_2[1728887:1725876]);
csa_3012 csau_3012_i789(tree_1[2596343:2593332],tree_1[2599355:2596344],tree_1[2602367:2599356],tree_2[1731899:1728888],tree_2[1734911:1731900]);
csa_3012 csau_3012_i790(tree_1[2605379:2602368],tree_1[2608391:2605380],tree_1[2611403:2608392],tree_2[1737923:1734912],tree_2[1740935:1737924]);
csa_3012 csau_3012_i791(tree_1[2614415:2611404],tree_1[2617427:2614416],tree_1[2620439:2617428],tree_2[1743947:1740936],tree_2[1746959:1743948]);
csa_3012 csau_3012_i792(tree_1[2623451:2620440],tree_1[2626463:2623452],tree_1[2629475:2626464],tree_2[1749971:1746960],tree_2[1752983:1749972]);
csa_3012 csau_3012_i793(tree_1[2632487:2629476],tree_1[2635499:2632488],tree_1[2638511:2635500],tree_2[1755995:1752984],tree_2[1759007:1755996]);
csa_3012 csau_3012_i794(tree_1[2641523:2638512],tree_1[2644535:2641524],tree_1[2647547:2644536],tree_2[1762019:1759008],tree_2[1765031:1762020]);
csa_3012 csau_3012_i795(tree_1[2650559:2647548],tree_1[2653571:2650560],tree_1[2656583:2653572],tree_2[1768043:1765032],tree_2[1771055:1768044]);
csa_3012 csau_3012_i796(tree_1[2659595:2656584],tree_1[2662607:2659596],tree_1[2665619:2662608],tree_2[1774067:1771056],tree_2[1777079:1774068]);
csa_3012 csau_3012_i797(tree_1[2668631:2665620],tree_1[2671643:2668632],tree_1[2674655:2671644],tree_2[1780091:1777080],tree_2[1783103:1780092]);
csa_3012 csau_3012_i798(tree_1[2677667:2674656],tree_1[2680679:2677668],tree_1[2683691:2680680],tree_2[1786115:1783104],tree_2[1789127:1786116]);
csa_3012 csau_3012_i799(tree_1[2686703:2683692],tree_1[2689715:2686704],tree_1[2692727:2689716],tree_2[1792139:1789128],tree_2[1795151:1792140]);
csa_3012 csau_3012_i800(tree_1[2695739:2692728],tree_1[2698751:2695740],tree_1[2701763:2698752],tree_2[1798163:1795152],tree_2[1801175:1798164]);
csa_3012 csau_3012_i801(tree_1[2704775:2701764],tree_1[2707787:2704776],tree_1[2710799:2707788],tree_2[1804187:1801176],tree_2[1807199:1804188]);
csa_3012 csau_3012_i802(tree_1[2713811:2710800],tree_1[2716823:2713812],tree_1[2719835:2716824],tree_2[1810211:1807200],tree_2[1813223:1810212]);
csa_3012 csau_3012_i803(tree_1[2722847:2719836],tree_1[2725859:2722848],tree_1[2728871:2725860],tree_2[1816235:1813224],tree_2[1819247:1816236]);
csa_3012 csau_3012_i804(tree_1[2731883:2728872],tree_1[2734895:2731884],tree_1[2737907:2734896],tree_2[1822259:1819248],tree_2[1825271:1822260]);
csa_3012 csau_3012_i805(tree_1[2740919:2737908],tree_1[2743931:2740920],tree_1[2746943:2743932],tree_2[1828283:1825272],tree_2[1831295:1828284]);
csa_3012 csau_3012_i806(tree_1[2749955:2746944],tree_1[2752967:2749956],tree_1[2755979:2752968],tree_2[1834307:1831296],tree_2[1837319:1834308]);
csa_3012 csau_3012_i807(tree_1[2758991:2755980],tree_1[2762003:2758992],tree_1[2765015:2762004],tree_2[1840331:1837320],tree_2[1843343:1840332]);
csa_3012 csau_3012_i808(tree_1[2768027:2765016],tree_1[2771039:2768028],tree_1[2774051:2771040],tree_2[1846355:1843344],tree_2[1849367:1846356]);
csa_3012 csau_3012_i809(tree_1[2777063:2774052],tree_1[2780075:2777064],tree_1[2783087:2780076],tree_2[1852379:1849368],tree_2[1855391:1852380]);
csa_3012 csau_3012_i810(tree_1[2786099:2783088],tree_1[2789111:2786100],tree_1[2792123:2789112],tree_2[1858403:1855392],tree_2[1861415:1858404]);
csa_3012 csau_3012_i811(tree_1[2795135:2792124],tree_1[2798147:2795136],tree_1[2801159:2798148],tree_2[1864427:1861416],tree_2[1867439:1864428]);
csa_3012 csau_3012_i812(tree_1[2804171:2801160],tree_1[2807183:2804172],tree_1[2810195:2807184],tree_2[1870451:1867440],tree_2[1873463:1870452]);
csa_3012 csau_3012_i813(tree_1[2813207:2810196],tree_1[2816219:2813208],tree_1[2819231:2816220],tree_2[1876475:1873464],tree_2[1879487:1876476]);
csa_3012 csau_3012_i814(tree_1[2822243:2819232],tree_1[2825255:2822244],tree_1[2828267:2825256],tree_2[1882499:1879488],tree_2[1885511:1882500]);
csa_3012 csau_3012_i815(tree_1[2831279:2828268],tree_1[2834291:2831280],tree_1[2837303:2834292],tree_2[1888523:1885512],tree_2[1891535:1888524]);
csa_3012 csau_3012_i816(tree_1[2840315:2837304],tree_1[2843327:2840316],tree_1[2846339:2843328],tree_2[1894547:1891536],tree_2[1897559:1894548]);
csa_3012 csau_3012_i817(tree_1[2849351:2846340],tree_1[2852363:2849352],tree_1[2855375:2852364],tree_2[1900571:1897560],tree_2[1903583:1900572]);
csa_3012 csau_3012_i818(tree_1[2858387:2855376],tree_1[2861399:2858388],tree_1[2864411:2861400],tree_2[1906595:1903584],tree_2[1909607:1906596]);
csa_3012 csau_3012_i819(tree_1[2867423:2864412],tree_1[2870435:2867424],tree_1[2873447:2870436],tree_2[1912619:1909608],tree_2[1915631:1912620]);
csa_3012 csau_3012_i820(tree_1[2876459:2873448],tree_1[2879471:2876460],tree_1[2882483:2879472],tree_2[1918643:1915632],tree_2[1921655:1918644]);
csa_3012 csau_3012_i821(tree_1[2885495:2882484],tree_1[2888507:2885496],tree_1[2891519:2888508],tree_2[1924667:1921656],tree_2[1927679:1924668]);
csa_3012 csau_3012_i822(tree_1[2894531:2891520],tree_1[2897543:2894532],tree_1[2900555:2897544],tree_2[1930691:1927680],tree_2[1933703:1930692]);
csa_3012 csau_3012_i823(tree_1[2903567:2900556],tree_1[2906579:2903568],tree_1[2909591:2906580],tree_2[1936715:1933704],tree_2[1939727:1936716]);
csa_3012 csau_3012_i824(tree_1[2912603:2909592],tree_1[2915615:2912604],tree_1[2918627:2915616],tree_2[1942739:1939728],tree_2[1945751:1942740]);
csa_3012 csau_3012_i825(tree_1[2921639:2918628],tree_1[2924651:2921640],tree_1[2927663:2924652],tree_2[1948763:1945752],tree_2[1951775:1948764]);
csa_3012 csau_3012_i826(tree_1[2930675:2927664],tree_1[2933687:2930676],tree_1[2936699:2933688],tree_2[1954787:1951776],tree_2[1957799:1954788]);
csa_3012 csau_3012_i827(tree_1[2939711:2936700],tree_1[2942723:2939712],tree_1[2945735:2942724],tree_2[1960811:1957800],tree_2[1963823:1960812]);
csa_3012 csau_3012_i828(tree_1[2948747:2945736],tree_1[2951759:2948748],tree_1[2954771:2951760],tree_2[1966835:1963824],tree_2[1969847:1966836]);
csa_3012 csau_3012_i829(tree_1[2957783:2954772],tree_1[2960795:2957784],tree_1[2963807:2960796],tree_2[1972859:1969848],tree_2[1975871:1972860]);
csa_3012 csau_3012_i830(tree_1[2966819:2963808],tree_1[2969831:2966820],tree_1[2972843:2969832],tree_2[1978883:1975872],tree_2[1981895:1978884]);
csa_3012 csau_3012_i831(tree_1[2975855:2972844],tree_1[2978867:2975856],tree_1[2981879:2978868],tree_2[1984907:1981896],tree_2[1987919:1984908]);
csa_3012 csau_3012_i832(tree_1[2984891:2981880],tree_1[2987903:2984892],tree_1[2990915:2987904],tree_2[1990931:1987920],tree_2[1993943:1990932]);
csa_3012 csau_3012_i833(tree_1[2993927:2990916],tree_1[2996939:2993928],tree_1[2999951:2996940],tree_2[1996955:1993944],tree_2[1999967:1996956]);
csa_3012 csau_3012_i834(tree_1[3002963:2999952],tree_1[3005975:3002964],tree_1[3008987:3005976],tree_2[2002979:1999968],tree_2[2005991:2002980]);
csa_3012 csau_3012_i835(tree_1[3011999:3008988],tree_1[3015011:3012000],tree_1[3018023:3015012],tree_2[2009003:2005992],tree_2[2012015:2009004]);
assign tree_2[2015027:2012016] = tree_1[3021035:3018024];
assign tree_2[2018039:2015028] = tree_1[3024047:3021036];
// layer-3
csa_3012 csau_3012_i836(tree_2[3011:0],tree_2[6023:3012],tree_2[9035:6024],tree_3[3011:0],tree_3[6023:3012]);
csa_3012 csau_3012_i837(tree_2[12047:9036],tree_2[15059:12048],tree_2[18071:15060],tree_3[9035:6024],tree_3[12047:9036]);
csa_3012 csau_3012_i838(tree_2[21083:18072],tree_2[24095:21084],tree_2[27107:24096],tree_3[15059:12048],tree_3[18071:15060]);
csa_3012 csau_3012_i839(tree_2[30119:27108],tree_2[33131:30120],tree_2[36143:33132],tree_3[21083:18072],tree_3[24095:21084]);
csa_3012 csau_3012_i840(tree_2[39155:36144],tree_2[42167:39156],tree_2[45179:42168],tree_3[27107:24096],tree_3[30119:27108]);
csa_3012 csau_3012_i841(tree_2[48191:45180],tree_2[51203:48192],tree_2[54215:51204],tree_3[33131:30120],tree_3[36143:33132]);
csa_3012 csau_3012_i842(tree_2[57227:54216],tree_2[60239:57228],tree_2[63251:60240],tree_3[39155:36144],tree_3[42167:39156]);
csa_3012 csau_3012_i843(tree_2[66263:63252],tree_2[69275:66264],tree_2[72287:69276],tree_3[45179:42168],tree_3[48191:45180]);
csa_3012 csau_3012_i844(tree_2[75299:72288],tree_2[78311:75300],tree_2[81323:78312],tree_3[51203:48192],tree_3[54215:51204]);
csa_3012 csau_3012_i845(tree_2[84335:81324],tree_2[87347:84336],tree_2[90359:87348],tree_3[57227:54216],tree_3[60239:57228]);
csa_3012 csau_3012_i846(tree_2[93371:90360],tree_2[96383:93372],tree_2[99395:96384],tree_3[63251:60240],tree_3[66263:63252]);
csa_3012 csau_3012_i847(tree_2[102407:99396],tree_2[105419:102408],tree_2[108431:105420],tree_3[69275:66264],tree_3[72287:69276]);
csa_3012 csau_3012_i848(tree_2[111443:108432],tree_2[114455:111444],tree_2[117467:114456],tree_3[75299:72288],tree_3[78311:75300]);
csa_3012 csau_3012_i849(tree_2[120479:117468],tree_2[123491:120480],tree_2[126503:123492],tree_3[81323:78312],tree_3[84335:81324]);
csa_3012 csau_3012_i850(tree_2[129515:126504],tree_2[132527:129516],tree_2[135539:132528],tree_3[87347:84336],tree_3[90359:87348]);
csa_3012 csau_3012_i851(tree_2[138551:135540],tree_2[141563:138552],tree_2[144575:141564],tree_3[93371:90360],tree_3[96383:93372]);
csa_3012 csau_3012_i852(tree_2[147587:144576],tree_2[150599:147588],tree_2[153611:150600],tree_3[99395:96384],tree_3[102407:99396]);
csa_3012 csau_3012_i853(tree_2[156623:153612],tree_2[159635:156624],tree_2[162647:159636],tree_3[105419:102408],tree_3[108431:105420]);
csa_3012 csau_3012_i854(tree_2[165659:162648],tree_2[168671:165660],tree_2[171683:168672],tree_3[111443:108432],tree_3[114455:111444]);
csa_3012 csau_3012_i855(tree_2[174695:171684],tree_2[177707:174696],tree_2[180719:177708],tree_3[117467:114456],tree_3[120479:117468]);
csa_3012 csau_3012_i856(tree_2[183731:180720],tree_2[186743:183732],tree_2[189755:186744],tree_3[123491:120480],tree_3[126503:123492]);
csa_3012 csau_3012_i857(tree_2[192767:189756],tree_2[195779:192768],tree_2[198791:195780],tree_3[129515:126504],tree_3[132527:129516]);
csa_3012 csau_3012_i858(tree_2[201803:198792],tree_2[204815:201804],tree_2[207827:204816],tree_3[135539:132528],tree_3[138551:135540]);
csa_3012 csau_3012_i859(tree_2[210839:207828],tree_2[213851:210840],tree_2[216863:213852],tree_3[141563:138552],tree_3[144575:141564]);
csa_3012 csau_3012_i860(tree_2[219875:216864],tree_2[222887:219876],tree_2[225899:222888],tree_3[147587:144576],tree_3[150599:147588]);
csa_3012 csau_3012_i861(tree_2[228911:225900],tree_2[231923:228912],tree_2[234935:231924],tree_3[153611:150600],tree_3[156623:153612]);
csa_3012 csau_3012_i862(tree_2[237947:234936],tree_2[240959:237948],tree_2[243971:240960],tree_3[159635:156624],tree_3[162647:159636]);
csa_3012 csau_3012_i863(tree_2[246983:243972],tree_2[249995:246984],tree_2[253007:249996],tree_3[165659:162648],tree_3[168671:165660]);
csa_3012 csau_3012_i864(tree_2[256019:253008],tree_2[259031:256020],tree_2[262043:259032],tree_3[171683:168672],tree_3[174695:171684]);
csa_3012 csau_3012_i865(tree_2[265055:262044],tree_2[268067:265056],tree_2[271079:268068],tree_3[177707:174696],tree_3[180719:177708]);
csa_3012 csau_3012_i866(tree_2[274091:271080],tree_2[277103:274092],tree_2[280115:277104],tree_3[183731:180720],tree_3[186743:183732]);
csa_3012 csau_3012_i867(tree_2[283127:280116],tree_2[286139:283128],tree_2[289151:286140],tree_3[189755:186744],tree_3[192767:189756]);
csa_3012 csau_3012_i868(tree_2[292163:289152],tree_2[295175:292164],tree_2[298187:295176],tree_3[195779:192768],tree_3[198791:195780]);
csa_3012 csau_3012_i869(tree_2[301199:298188],tree_2[304211:301200],tree_2[307223:304212],tree_3[201803:198792],tree_3[204815:201804]);
csa_3012 csau_3012_i870(tree_2[310235:307224],tree_2[313247:310236],tree_2[316259:313248],tree_3[207827:204816],tree_3[210839:207828]);
csa_3012 csau_3012_i871(tree_2[319271:316260],tree_2[322283:319272],tree_2[325295:322284],tree_3[213851:210840],tree_3[216863:213852]);
csa_3012 csau_3012_i872(tree_2[328307:325296],tree_2[331319:328308],tree_2[334331:331320],tree_3[219875:216864],tree_3[222887:219876]);
csa_3012 csau_3012_i873(tree_2[337343:334332],tree_2[340355:337344],tree_2[343367:340356],tree_3[225899:222888],tree_3[228911:225900]);
csa_3012 csau_3012_i874(tree_2[346379:343368],tree_2[349391:346380],tree_2[352403:349392],tree_3[231923:228912],tree_3[234935:231924]);
csa_3012 csau_3012_i875(tree_2[355415:352404],tree_2[358427:355416],tree_2[361439:358428],tree_3[237947:234936],tree_3[240959:237948]);
csa_3012 csau_3012_i876(tree_2[364451:361440],tree_2[367463:364452],tree_2[370475:367464],tree_3[243971:240960],tree_3[246983:243972]);
csa_3012 csau_3012_i877(tree_2[373487:370476],tree_2[376499:373488],tree_2[379511:376500],tree_3[249995:246984],tree_3[253007:249996]);
csa_3012 csau_3012_i878(tree_2[382523:379512],tree_2[385535:382524],tree_2[388547:385536],tree_3[256019:253008],tree_3[259031:256020]);
csa_3012 csau_3012_i879(tree_2[391559:388548],tree_2[394571:391560],tree_2[397583:394572],tree_3[262043:259032],tree_3[265055:262044]);
csa_3012 csau_3012_i880(tree_2[400595:397584],tree_2[403607:400596],tree_2[406619:403608],tree_3[268067:265056],tree_3[271079:268068]);
csa_3012 csau_3012_i881(tree_2[409631:406620],tree_2[412643:409632],tree_2[415655:412644],tree_3[274091:271080],tree_3[277103:274092]);
csa_3012 csau_3012_i882(tree_2[418667:415656],tree_2[421679:418668],tree_2[424691:421680],tree_3[280115:277104],tree_3[283127:280116]);
csa_3012 csau_3012_i883(tree_2[427703:424692],tree_2[430715:427704],tree_2[433727:430716],tree_3[286139:283128],tree_3[289151:286140]);
csa_3012 csau_3012_i884(tree_2[436739:433728],tree_2[439751:436740],tree_2[442763:439752],tree_3[292163:289152],tree_3[295175:292164]);
csa_3012 csau_3012_i885(tree_2[445775:442764],tree_2[448787:445776],tree_2[451799:448788],tree_3[298187:295176],tree_3[301199:298188]);
csa_3012 csau_3012_i886(tree_2[454811:451800],tree_2[457823:454812],tree_2[460835:457824],tree_3[304211:301200],tree_3[307223:304212]);
csa_3012 csau_3012_i887(tree_2[463847:460836],tree_2[466859:463848],tree_2[469871:466860],tree_3[310235:307224],tree_3[313247:310236]);
csa_3012 csau_3012_i888(tree_2[472883:469872],tree_2[475895:472884],tree_2[478907:475896],tree_3[316259:313248],tree_3[319271:316260]);
csa_3012 csau_3012_i889(tree_2[481919:478908],tree_2[484931:481920],tree_2[487943:484932],tree_3[322283:319272],tree_3[325295:322284]);
csa_3012 csau_3012_i890(tree_2[490955:487944],tree_2[493967:490956],tree_2[496979:493968],tree_3[328307:325296],tree_3[331319:328308]);
csa_3012 csau_3012_i891(tree_2[499991:496980],tree_2[503003:499992],tree_2[506015:503004],tree_3[334331:331320],tree_3[337343:334332]);
csa_3012 csau_3012_i892(tree_2[509027:506016],tree_2[512039:509028],tree_2[515051:512040],tree_3[340355:337344],tree_3[343367:340356]);
csa_3012 csau_3012_i893(tree_2[518063:515052],tree_2[521075:518064],tree_2[524087:521076],tree_3[346379:343368],tree_3[349391:346380]);
csa_3012 csau_3012_i894(tree_2[527099:524088],tree_2[530111:527100],tree_2[533123:530112],tree_3[352403:349392],tree_3[355415:352404]);
csa_3012 csau_3012_i895(tree_2[536135:533124],tree_2[539147:536136],tree_2[542159:539148],tree_3[358427:355416],tree_3[361439:358428]);
csa_3012 csau_3012_i896(tree_2[545171:542160],tree_2[548183:545172],tree_2[551195:548184],tree_3[364451:361440],tree_3[367463:364452]);
csa_3012 csau_3012_i897(tree_2[554207:551196],tree_2[557219:554208],tree_2[560231:557220],tree_3[370475:367464],tree_3[373487:370476]);
csa_3012 csau_3012_i898(tree_2[563243:560232],tree_2[566255:563244],tree_2[569267:566256],tree_3[376499:373488],tree_3[379511:376500]);
csa_3012 csau_3012_i899(tree_2[572279:569268],tree_2[575291:572280],tree_2[578303:575292],tree_3[382523:379512],tree_3[385535:382524]);
csa_3012 csau_3012_i900(tree_2[581315:578304],tree_2[584327:581316],tree_2[587339:584328],tree_3[388547:385536],tree_3[391559:388548]);
csa_3012 csau_3012_i901(tree_2[590351:587340],tree_2[593363:590352],tree_2[596375:593364],tree_3[394571:391560],tree_3[397583:394572]);
csa_3012 csau_3012_i902(tree_2[599387:596376],tree_2[602399:599388],tree_2[605411:602400],tree_3[400595:397584],tree_3[403607:400596]);
csa_3012 csau_3012_i903(tree_2[608423:605412],tree_2[611435:608424],tree_2[614447:611436],tree_3[406619:403608],tree_3[409631:406620]);
csa_3012 csau_3012_i904(tree_2[617459:614448],tree_2[620471:617460],tree_2[623483:620472],tree_3[412643:409632],tree_3[415655:412644]);
csa_3012 csau_3012_i905(tree_2[626495:623484],tree_2[629507:626496],tree_2[632519:629508],tree_3[418667:415656],tree_3[421679:418668]);
csa_3012 csau_3012_i906(tree_2[635531:632520],tree_2[638543:635532],tree_2[641555:638544],tree_3[424691:421680],tree_3[427703:424692]);
csa_3012 csau_3012_i907(tree_2[644567:641556],tree_2[647579:644568],tree_2[650591:647580],tree_3[430715:427704],tree_3[433727:430716]);
csa_3012 csau_3012_i908(tree_2[653603:650592],tree_2[656615:653604],tree_2[659627:656616],tree_3[436739:433728],tree_3[439751:436740]);
csa_3012 csau_3012_i909(tree_2[662639:659628],tree_2[665651:662640],tree_2[668663:665652],tree_3[442763:439752],tree_3[445775:442764]);
csa_3012 csau_3012_i910(tree_2[671675:668664],tree_2[674687:671676],tree_2[677699:674688],tree_3[448787:445776],tree_3[451799:448788]);
csa_3012 csau_3012_i911(tree_2[680711:677700],tree_2[683723:680712],tree_2[686735:683724],tree_3[454811:451800],tree_3[457823:454812]);
csa_3012 csau_3012_i912(tree_2[689747:686736],tree_2[692759:689748],tree_2[695771:692760],tree_3[460835:457824],tree_3[463847:460836]);
csa_3012 csau_3012_i913(tree_2[698783:695772],tree_2[701795:698784],tree_2[704807:701796],tree_3[466859:463848],tree_3[469871:466860]);
csa_3012 csau_3012_i914(tree_2[707819:704808],tree_2[710831:707820],tree_2[713843:710832],tree_3[472883:469872],tree_3[475895:472884]);
csa_3012 csau_3012_i915(tree_2[716855:713844],tree_2[719867:716856],tree_2[722879:719868],tree_3[478907:475896],tree_3[481919:478908]);
csa_3012 csau_3012_i916(tree_2[725891:722880],tree_2[728903:725892],tree_2[731915:728904],tree_3[484931:481920],tree_3[487943:484932]);
csa_3012 csau_3012_i917(tree_2[734927:731916],tree_2[737939:734928],tree_2[740951:737940],tree_3[490955:487944],tree_3[493967:490956]);
csa_3012 csau_3012_i918(tree_2[743963:740952],tree_2[746975:743964],tree_2[749987:746976],tree_3[496979:493968],tree_3[499991:496980]);
csa_3012 csau_3012_i919(tree_2[752999:749988],tree_2[756011:753000],tree_2[759023:756012],tree_3[503003:499992],tree_3[506015:503004]);
csa_3012 csau_3012_i920(tree_2[762035:759024],tree_2[765047:762036],tree_2[768059:765048],tree_3[509027:506016],tree_3[512039:509028]);
csa_3012 csau_3012_i921(tree_2[771071:768060],tree_2[774083:771072],tree_2[777095:774084],tree_3[515051:512040],tree_3[518063:515052]);
csa_3012 csau_3012_i922(tree_2[780107:777096],tree_2[783119:780108],tree_2[786131:783120],tree_3[521075:518064],tree_3[524087:521076]);
csa_3012 csau_3012_i923(tree_2[789143:786132],tree_2[792155:789144],tree_2[795167:792156],tree_3[527099:524088],tree_3[530111:527100]);
csa_3012 csau_3012_i924(tree_2[798179:795168],tree_2[801191:798180],tree_2[804203:801192],tree_3[533123:530112],tree_3[536135:533124]);
csa_3012 csau_3012_i925(tree_2[807215:804204],tree_2[810227:807216],tree_2[813239:810228],tree_3[539147:536136],tree_3[542159:539148]);
csa_3012 csau_3012_i926(tree_2[816251:813240],tree_2[819263:816252],tree_2[822275:819264],tree_3[545171:542160],tree_3[548183:545172]);
csa_3012 csau_3012_i927(tree_2[825287:822276],tree_2[828299:825288],tree_2[831311:828300],tree_3[551195:548184],tree_3[554207:551196]);
csa_3012 csau_3012_i928(tree_2[834323:831312],tree_2[837335:834324],tree_2[840347:837336],tree_3[557219:554208],tree_3[560231:557220]);
csa_3012 csau_3012_i929(tree_2[843359:840348],tree_2[846371:843360],tree_2[849383:846372],tree_3[563243:560232],tree_3[566255:563244]);
csa_3012 csau_3012_i930(tree_2[852395:849384],tree_2[855407:852396],tree_2[858419:855408],tree_3[569267:566256],tree_3[572279:569268]);
csa_3012 csau_3012_i931(tree_2[861431:858420],tree_2[864443:861432],tree_2[867455:864444],tree_3[575291:572280],tree_3[578303:575292]);
csa_3012 csau_3012_i932(tree_2[870467:867456],tree_2[873479:870468],tree_2[876491:873480],tree_3[581315:578304],tree_3[584327:581316]);
csa_3012 csau_3012_i933(tree_2[879503:876492],tree_2[882515:879504],tree_2[885527:882516],tree_3[587339:584328],tree_3[590351:587340]);
csa_3012 csau_3012_i934(tree_2[888539:885528],tree_2[891551:888540],tree_2[894563:891552],tree_3[593363:590352],tree_3[596375:593364]);
csa_3012 csau_3012_i935(tree_2[897575:894564],tree_2[900587:897576],tree_2[903599:900588],tree_3[599387:596376],tree_3[602399:599388]);
csa_3012 csau_3012_i936(tree_2[906611:903600],tree_2[909623:906612],tree_2[912635:909624],tree_3[605411:602400],tree_3[608423:605412]);
csa_3012 csau_3012_i937(tree_2[915647:912636],tree_2[918659:915648],tree_2[921671:918660],tree_3[611435:608424],tree_3[614447:611436]);
csa_3012 csau_3012_i938(tree_2[924683:921672],tree_2[927695:924684],tree_2[930707:927696],tree_3[617459:614448],tree_3[620471:617460]);
csa_3012 csau_3012_i939(tree_2[933719:930708],tree_2[936731:933720],tree_2[939743:936732],tree_3[623483:620472],tree_3[626495:623484]);
csa_3012 csau_3012_i940(tree_2[942755:939744],tree_2[945767:942756],tree_2[948779:945768],tree_3[629507:626496],tree_3[632519:629508]);
csa_3012 csau_3012_i941(tree_2[951791:948780],tree_2[954803:951792],tree_2[957815:954804],tree_3[635531:632520],tree_3[638543:635532]);
csa_3012 csau_3012_i942(tree_2[960827:957816],tree_2[963839:960828],tree_2[966851:963840],tree_3[641555:638544],tree_3[644567:641556]);
csa_3012 csau_3012_i943(tree_2[969863:966852],tree_2[972875:969864],tree_2[975887:972876],tree_3[647579:644568],tree_3[650591:647580]);
csa_3012 csau_3012_i944(tree_2[978899:975888],tree_2[981911:978900],tree_2[984923:981912],tree_3[653603:650592],tree_3[656615:653604]);
csa_3012 csau_3012_i945(tree_2[987935:984924],tree_2[990947:987936],tree_2[993959:990948],tree_3[659627:656616],tree_3[662639:659628]);
csa_3012 csau_3012_i946(tree_2[996971:993960],tree_2[999983:996972],tree_2[1002995:999984],tree_3[665651:662640],tree_3[668663:665652]);
csa_3012 csau_3012_i947(tree_2[1006007:1002996],tree_2[1009019:1006008],tree_2[1012031:1009020],tree_3[671675:668664],tree_3[674687:671676]);
csa_3012 csau_3012_i948(tree_2[1015043:1012032],tree_2[1018055:1015044],tree_2[1021067:1018056],tree_3[677699:674688],tree_3[680711:677700]);
csa_3012 csau_3012_i949(tree_2[1024079:1021068],tree_2[1027091:1024080],tree_2[1030103:1027092],tree_3[683723:680712],tree_3[686735:683724]);
csa_3012 csau_3012_i950(tree_2[1033115:1030104],tree_2[1036127:1033116],tree_2[1039139:1036128],tree_3[689747:686736],tree_3[692759:689748]);
csa_3012 csau_3012_i951(tree_2[1042151:1039140],tree_2[1045163:1042152],tree_2[1048175:1045164],tree_3[695771:692760],tree_3[698783:695772]);
csa_3012 csau_3012_i952(tree_2[1051187:1048176],tree_2[1054199:1051188],tree_2[1057211:1054200],tree_3[701795:698784],tree_3[704807:701796]);
csa_3012 csau_3012_i953(tree_2[1060223:1057212],tree_2[1063235:1060224],tree_2[1066247:1063236],tree_3[707819:704808],tree_3[710831:707820]);
csa_3012 csau_3012_i954(tree_2[1069259:1066248],tree_2[1072271:1069260],tree_2[1075283:1072272],tree_3[713843:710832],tree_3[716855:713844]);
csa_3012 csau_3012_i955(tree_2[1078295:1075284],tree_2[1081307:1078296],tree_2[1084319:1081308],tree_3[719867:716856],tree_3[722879:719868]);
csa_3012 csau_3012_i956(tree_2[1087331:1084320],tree_2[1090343:1087332],tree_2[1093355:1090344],tree_3[725891:722880],tree_3[728903:725892]);
csa_3012 csau_3012_i957(tree_2[1096367:1093356],tree_2[1099379:1096368],tree_2[1102391:1099380],tree_3[731915:728904],tree_3[734927:731916]);
csa_3012 csau_3012_i958(tree_2[1105403:1102392],tree_2[1108415:1105404],tree_2[1111427:1108416],tree_3[737939:734928],tree_3[740951:737940]);
csa_3012 csau_3012_i959(tree_2[1114439:1111428],tree_2[1117451:1114440],tree_2[1120463:1117452],tree_3[743963:740952],tree_3[746975:743964]);
csa_3012 csau_3012_i960(tree_2[1123475:1120464],tree_2[1126487:1123476],tree_2[1129499:1126488],tree_3[749987:746976],tree_3[752999:749988]);
csa_3012 csau_3012_i961(tree_2[1132511:1129500],tree_2[1135523:1132512],tree_2[1138535:1135524],tree_3[756011:753000],tree_3[759023:756012]);
csa_3012 csau_3012_i962(tree_2[1141547:1138536],tree_2[1144559:1141548],tree_2[1147571:1144560],tree_3[762035:759024],tree_3[765047:762036]);
csa_3012 csau_3012_i963(tree_2[1150583:1147572],tree_2[1153595:1150584],tree_2[1156607:1153596],tree_3[768059:765048],tree_3[771071:768060]);
csa_3012 csau_3012_i964(tree_2[1159619:1156608],tree_2[1162631:1159620],tree_2[1165643:1162632],tree_3[774083:771072],tree_3[777095:774084]);
csa_3012 csau_3012_i965(tree_2[1168655:1165644],tree_2[1171667:1168656],tree_2[1174679:1171668],tree_3[780107:777096],tree_3[783119:780108]);
csa_3012 csau_3012_i966(tree_2[1177691:1174680],tree_2[1180703:1177692],tree_2[1183715:1180704],tree_3[786131:783120],tree_3[789143:786132]);
csa_3012 csau_3012_i967(tree_2[1186727:1183716],tree_2[1189739:1186728],tree_2[1192751:1189740],tree_3[792155:789144],tree_3[795167:792156]);
csa_3012 csau_3012_i968(tree_2[1195763:1192752],tree_2[1198775:1195764],tree_2[1201787:1198776],tree_3[798179:795168],tree_3[801191:798180]);
csa_3012 csau_3012_i969(tree_2[1204799:1201788],tree_2[1207811:1204800],tree_2[1210823:1207812],tree_3[804203:801192],tree_3[807215:804204]);
csa_3012 csau_3012_i970(tree_2[1213835:1210824],tree_2[1216847:1213836],tree_2[1219859:1216848],tree_3[810227:807216],tree_3[813239:810228]);
csa_3012 csau_3012_i971(tree_2[1222871:1219860],tree_2[1225883:1222872],tree_2[1228895:1225884],tree_3[816251:813240],tree_3[819263:816252]);
csa_3012 csau_3012_i972(tree_2[1231907:1228896],tree_2[1234919:1231908],tree_2[1237931:1234920],tree_3[822275:819264],tree_3[825287:822276]);
csa_3012 csau_3012_i973(tree_2[1240943:1237932],tree_2[1243955:1240944],tree_2[1246967:1243956],tree_3[828299:825288],tree_3[831311:828300]);
csa_3012 csau_3012_i974(tree_2[1249979:1246968],tree_2[1252991:1249980],tree_2[1256003:1252992],tree_3[834323:831312],tree_3[837335:834324]);
csa_3012 csau_3012_i975(tree_2[1259015:1256004],tree_2[1262027:1259016],tree_2[1265039:1262028],tree_3[840347:837336],tree_3[843359:840348]);
csa_3012 csau_3012_i976(tree_2[1268051:1265040],tree_2[1271063:1268052],tree_2[1274075:1271064],tree_3[846371:843360],tree_3[849383:846372]);
csa_3012 csau_3012_i977(tree_2[1277087:1274076],tree_2[1280099:1277088],tree_2[1283111:1280100],tree_3[852395:849384],tree_3[855407:852396]);
csa_3012 csau_3012_i978(tree_2[1286123:1283112],tree_2[1289135:1286124],tree_2[1292147:1289136],tree_3[858419:855408],tree_3[861431:858420]);
csa_3012 csau_3012_i979(tree_2[1295159:1292148],tree_2[1298171:1295160],tree_2[1301183:1298172],tree_3[864443:861432],tree_3[867455:864444]);
csa_3012 csau_3012_i980(tree_2[1304195:1301184],tree_2[1307207:1304196],tree_2[1310219:1307208],tree_3[870467:867456],tree_3[873479:870468]);
csa_3012 csau_3012_i981(tree_2[1313231:1310220],tree_2[1316243:1313232],tree_2[1319255:1316244],tree_3[876491:873480],tree_3[879503:876492]);
csa_3012 csau_3012_i982(tree_2[1322267:1319256],tree_2[1325279:1322268],tree_2[1328291:1325280],tree_3[882515:879504],tree_3[885527:882516]);
csa_3012 csau_3012_i983(tree_2[1331303:1328292],tree_2[1334315:1331304],tree_2[1337327:1334316],tree_3[888539:885528],tree_3[891551:888540]);
csa_3012 csau_3012_i984(tree_2[1340339:1337328],tree_2[1343351:1340340],tree_2[1346363:1343352],tree_3[894563:891552],tree_3[897575:894564]);
csa_3012 csau_3012_i985(tree_2[1349375:1346364],tree_2[1352387:1349376],tree_2[1355399:1352388],tree_3[900587:897576],tree_3[903599:900588]);
csa_3012 csau_3012_i986(tree_2[1358411:1355400],tree_2[1361423:1358412],tree_2[1364435:1361424],tree_3[906611:903600],tree_3[909623:906612]);
csa_3012 csau_3012_i987(tree_2[1367447:1364436],tree_2[1370459:1367448],tree_2[1373471:1370460],tree_3[912635:909624],tree_3[915647:912636]);
csa_3012 csau_3012_i988(tree_2[1376483:1373472],tree_2[1379495:1376484],tree_2[1382507:1379496],tree_3[918659:915648],tree_3[921671:918660]);
csa_3012 csau_3012_i989(tree_2[1385519:1382508],tree_2[1388531:1385520],tree_2[1391543:1388532],tree_3[924683:921672],tree_3[927695:924684]);
csa_3012 csau_3012_i990(tree_2[1394555:1391544],tree_2[1397567:1394556],tree_2[1400579:1397568],tree_3[930707:927696],tree_3[933719:930708]);
csa_3012 csau_3012_i991(tree_2[1403591:1400580],tree_2[1406603:1403592],tree_2[1409615:1406604],tree_3[936731:933720],tree_3[939743:936732]);
csa_3012 csau_3012_i992(tree_2[1412627:1409616],tree_2[1415639:1412628],tree_2[1418651:1415640],tree_3[942755:939744],tree_3[945767:942756]);
csa_3012 csau_3012_i993(tree_2[1421663:1418652],tree_2[1424675:1421664],tree_2[1427687:1424676],tree_3[948779:945768],tree_3[951791:948780]);
csa_3012 csau_3012_i994(tree_2[1430699:1427688],tree_2[1433711:1430700],tree_2[1436723:1433712],tree_3[954803:951792],tree_3[957815:954804]);
csa_3012 csau_3012_i995(tree_2[1439735:1436724],tree_2[1442747:1439736],tree_2[1445759:1442748],tree_3[960827:957816],tree_3[963839:960828]);
csa_3012 csau_3012_i996(tree_2[1448771:1445760],tree_2[1451783:1448772],tree_2[1454795:1451784],tree_3[966851:963840],tree_3[969863:966852]);
csa_3012 csau_3012_i997(tree_2[1457807:1454796],tree_2[1460819:1457808],tree_2[1463831:1460820],tree_3[972875:969864],tree_3[975887:972876]);
csa_3012 csau_3012_i998(tree_2[1466843:1463832],tree_2[1469855:1466844],tree_2[1472867:1469856],tree_3[978899:975888],tree_3[981911:978900]);
csa_3012 csau_3012_i999(tree_2[1475879:1472868],tree_2[1478891:1475880],tree_2[1481903:1478892],tree_3[984923:981912],tree_3[987935:984924]);
csa_3012 csau_3012_i1000(tree_2[1484915:1481904],tree_2[1487927:1484916],tree_2[1490939:1487928],tree_3[990947:987936],tree_3[993959:990948]);
csa_3012 csau_3012_i1001(tree_2[1493951:1490940],tree_2[1496963:1493952],tree_2[1499975:1496964],tree_3[996971:993960],tree_3[999983:996972]);
csa_3012 csau_3012_i1002(tree_2[1502987:1499976],tree_2[1505999:1502988],tree_2[1509011:1506000],tree_3[1002995:999984],tree_3[1006007:1002996]);
csa_3012 csau_3012_i1003(tree_2[1512023:1509012],tree_2[1515035:1512024],tree_2[1518047:1515036],tree_3[1009019:1006008],tree_3[1012031:1009020]);
csa_3012 csau_3012_i1004(tree_2[1521059:1518048],tree_2[1524071:1521060],tree_2[1527083:1524072],tree_3[1015043:1012032],tree_3[1018055:1015044]);
csa_3012 csau_3012_i1005(tree_2[1530095:1527084],tree_2[1533107:1530096],tree_2[1536119:1533108],tree_3[1021067:1018056],tree_3[1024079:1021068]);
csa_3012 csau_3012_i1006(tree_2[1539131:1536120],tree_2[1542143:1539132],tree_2[1545155:1542144],tree_3[1027091:1024080],tree_3[1030103:1027092]);
csa_3012 csau_3012_i1007(tree_2[1548167:1545156],tree_2[1551179:1548168],tree_2[1554191:1551180],tree_3[1033115:1030104],tree_3[1036127:1033116]);
csa_3012 csau_3012_i1008(tree_2[1557203:1554192],tree_2[1560215:1557204],tree_2[1563227:1560216],tree_3[1039139:1036128],tree_3[1042151:1039140]);
csa_3012 csau_3012_i1009(tree_2[1566239:1563228],tree_2[1569251:1566240],tree_2[1572263:1569252],tree_3[1045163:1042152],tree_3[1048175:1045164]);
csa_3012 csau_3012_i1010(tree_2[1575275:1572264],tree_2[1578287:1575276],tree_2[1581299:1578288],tree_3[1051187:1048176],tree_3[1054199:1051188]);
csa_3012 csau_3012_i1011(tree_2[1584311:1581300],tree_2[1587323:1584312],tree_2[1590335:1587324],tree_3[1057211:1054200],tree_3[1060223:1057212]);
csa_3012 csau_3012_i1012(tree_2[1593347:1590336],tree_2[1596359:1593348],tree_2[1599371:1596360],tree_3[1063235:1060224],tree_3[1066247:1063236]);
csa_3012 csau_3012_i1013(tree_2[1602383:1599372],tree_2[1605395:1602384],tree_2[1608407:1605396],tree_3[1069259:1066248],tree_3[1072271:1069260]);
csa_3012 csau_3012_i1014(tree_2[1611419:1608408],tree_2[1614431:1611420],tree_2[1617443:1614432],tree_3[1075283:1072272],tree_3[1078295:1075284]);
csa_3012 csau_3012_i1015(tree_2[1620455:1617444],tree_2[1623467:1620456],tree_2[1626479:1623468],tree_3[1081307:1078296],tree_3[1084319:1081308]);
csa_3012 csau_3012_i1016(tree_2[1629491:1626480],tree_2[1632503:1629492],tree_2[1635515:1632504],tree_3[1087331:1084320],tree_3[1090343:1087332]);
csa_3012 csau_3012_i1017(tree_2[1638527:1635516],tree_2[1641539:1638528],tree_2[1644551:1641540],tree_3[1093355:1090344],tree_3[1096367:1093356]);
csa_3012 csau_3012_i1018(tree_2[1647563:1644552],tree_2[1650575:1647564],tree_2[1653587:1650576],tree_3[1099379:1096368],tree_3[1102391:1099380]);
csa_3012 csau_3012_i1019(tree_2[1656599:1653588],tree_2[1659611:1656600],tree_2[1662623:1659612],tree_3[1105403:1102392],tree_3[1108415:1105404]);
csa_3012 csau_3012_i1020(tree_2[1665635:1662624],tree_2[1668647:1665636],tree_2[1671659:1668648],tree_3[1111427:1108416],tree_3[1114439:1111428]);
csa_3012 csau_3012_i1021(tree_2[1674671:1671660],tree_2[1677683:1674672],tree_2[1680695:1677684],tree_3[1117451:1114440],tree_3[1120463:1117452]);
csa_3012 csau_3012_i1022(tree_2[1683707:1680696],tree_2[1686719:1683708],tree_2[1689731:1686720],tree_3[1123475:1120464],tree_3[1126487:1123476]);
csa_3012 csau_3012_i1023(tree_2[1692743:1689732],tree_2[1695755:1692744],tree_2[1698767:1695756],tree_3[1129499:1126488],tree_3[1132511:1129500]);
csa_3012 csau_3012_i1024(tree_2[1701779:1698768],tree_2[1704791:1701780],tree_2[1707803:1704792],tree_3[1135523:1132512],tree_3[1138535:1135524]);
csa_3012 csau_3012_i1025(tree_2[1710815:1707804],tree_2[1713827:1710816],tree_2[1716839:1713828],tree_3[1141547:1138536],tree_3[1144559:1141548]);
csa_3012 csau_3012_i1026(tree_2[1719851:1716840],tree_2[1722863:1719852],tree_2[1725875:1722864],tree_3[1147571:1144560],tree_3[1150583:1147572]);
csa_3012 csau_3012_i1027(tree_2[1728887:1725876],tree_2[1731899:1728888],tree_2[1734911:1731900],tree_3[1153595:1150584],tree_3[1156607:1153596]);
csa_3012 csau_3012_i1028(tree_2[1737923:1734912],tree_2[1740935:1737924],tree_2[1743947:1740936],tree_3[1159619:1156608],tree_3[1162631:1159620]);
csa_3012 csau_3012_i1029(tree_2[1746959:1743948],tree_2[1749971:1746960],tree_2[1752983:1749972],tree_3[1165643:1162632],tree_3[1168655:1165644]);
csa_3012 csau_3012_i1030(tree_2[1755995:1752984],tree_2[1759007:1755996],tree_2[1762019:1759008],tree_3[1171667:1168656],tree_3[1174679:1171668]);
csa_3012 csau_3012_i1031(tree_2[1765031:1762020],tree_2[1768043:1765032],tree_2[1771055:1768044],tree_3[1177691:1174680],tree_3[1180703:1177692]);
csa_3012 csau_3012_i1032(tree_2[1774067:1771056],tree_2[1777079:1774068],tree_2[1780091:1777080],tree_3[1183715:1180704],tree_3[1186727:1183716]);
csa_3012 csau_3012_i1033(tree_2[1783103:1780092],tree_2[1786115:1783104],tree_2[1789127:1786116],tree_3[1189739:1186728],tree_3[1192751:1189740]);
csa_3012 csau_3012_i1034(tree_2[1792139:1789128],tree_2[1795151:1792140],tree_2[1798163:1795152],tree_3[1195763:1192752],tree_3[1198775:1195764]);
csa_3012 csau_3012_i1035(tree_2[1801175:1798164],tree_2[1804187:1801176],tree_2[1807199:1804188],tree_3[1201787:1198776],tree_3[1204799:1201788]);
csa_3012 csau_3012_i1036(tree_2[1810211:1807200],tree_2[1813223:1810212],tree_2[1816235:1813224],tree_3[1207811:1204800],tree_3[1210823:1207812]);
csa_3012 csau_3012_i1037(tree_2[1819247:1816236],tree_2[1822259:1819248],tree_2[1825271:1822260],tree_3[1213835:1210824],tree_3[1216847:1213836]);
csa_3012 csau_3012_i1038(tree_2[1828283:1825272],tree_2[1831295:1828284],tree_2[1834307:1831296],tree_3[1219859:1216848],tree_3[1222871:1219860]);
csa_3012 csau_3012_i1039(tree_2[1837319:1834308],tree_2[1840331:1837320],tree_2[1843343:1840332],tree_3[1225883:1222872],tree_3[1228895:1225884]);
csa_3012 csau_3012_i1040(tree_2[1846355:1843344],tree_2[1849367:1846356],tree_2[1852379:1849368],tree_3[1231907:1228896],tree_3[1234919:1231908]);
csa_3012 csau_3012_i1041(tree_2[1855391:1852380],tree_2[1858403:1855392],tree_2[1861415:1858404],tree_3[1237931:1234920],tree_3[1240943:1237932]);
csa_3012 csau_3012_i1042(tree_2[1864427:1861416],tree_2[1867439:1864428],tree_2[1870451:1867440],tree_3[1243955:1240944],tree_3[1246967:1243956]);
csa_3012 csau_3012_i1043(tree_2[1873463:1870452],tree_2[1876475:1873464],tree_2[1879487:1876476],tree_3[1249979:1246968],tree_3[1252991:1249980]);
csa_3012 csau_3012_i1044(tree_2[1882499:1879488],tree_2[1885511:1882500],tree_2[1888523:1885512],tree_3[1256003:1252992],tree_3[1259015:1256004]);
csa_3012 csau_3012_i1045(tree_2[1891535:1888524],tree_2[1894547:1891536],tree_2[1897559:1894548],tree_3[1262027:1259016],tree_3[1265039:1262028]);
csa_3012 csau_3012_i1046(tree_2[1900571:1897560],tree_2[1903583:1900572],tree_2[1906595:1903584],tree_3[1268051:1265040],tree_3[1271063:1268052]);
csa_3012 csau_3012_i1047(tree_2[1909607:1906596],tree_2[1912619:1909608],tree_2[1915631:1912620],tree_3[1274075:1271064],tree_3[1277087:1274076]);
csa_3012 csau_3012_i1048(tree_2[1918643:1915632],tree_2[1921655:1918644],tree_2[1924667:1921656],tree_3[1280099:1277088],tree_3[1283111:1280100]);
csa_3012 csau_3012_i1049(tree_2[1927679:1924668],tree_2[1930691:1927680],tree_2[1933703:1930692],tree_3[1286123:1283112],tree_3[1289135:1286124]);
csa_3012 csau_3012_i1050(tree_2[1936715:1933704],tree_2[1939727:1936716],tree_2[1942739:1939728],tree_3[1292147:1289136],tree_3[1295159:1292148]);
csa_3012 csau_3012_i1051(tree_2[1945751:1942740],tree_2[1948763:1945752],tree_2[1951775:1948764],tree_3[1298171:1295160],tree_3[1301183:1298172]);
csa_3012 csau_3012_i1052(tree_2[1954787:1951776],tree_2[1957799:1954788],tree_2[1960811:1957800],tree_3[1304195:1301184],tree_3[1307207:1304196]);
csa_3012 csau_3012_i1053(tree_2[1963823:1960812],tree_2[1966835:1963824],tree_2[1969847:1966836],tree_3[1310219:1307208],tree_3[1313231:1310220]);
csa_3012 csau_3012_i1054(tree_2[1972859:1969848],tree_2[1975871:1972860],tree_2[1978883:1975872],tree_3[1316243:1313232],tree_3[1319255:1316244]);
csa_3012 csau_3012_i1055(tree_2[1981895:1978884],tree_2[1984907:1981896],tree_2[1987919:1984908],tree_3[1322267:1319256],tree_3[1325279:1322268]);
csa_3012 csau_3012_i1056(tree_2[1990931:1987920],tree_2[1993943:1990932],tree_2[1996955:1993944],tree_3[1328291:1325280],tree_3[1331303:1328292]);
csa_3012 csau_3012_i1057(tree_2[1999967:1996956],tree_2[2002979:1999968],tree_2[2005991:2002980],tree_3[1334315:1331304],tree_3[1337327:1334316]);
csa_3012 csau_3012_i1058(tree_2[2009003:2005992],tree_2[2012015:2009004],tree_2[2015027:2012016],tree_3[1340339:1337328],tree_3[1343351:1340340]);
assign tree_3[1346363:1343352] = tree_2[2018039:2015028];
// layer-4
csa_3012 csau_3012_i1059(tree_3[3011:0],tree_3[6023:3012],tree_3[9035:6024],tree_4[3011:0],tree_4[6023:3012]);
csa_3012 csau_3012_i1060(tree_3[12047:9036],tree_3[15059:12048],tree_3[18071:15060],tree_4[9035:6024],tree_4[12047:9036]);
csa_3012 csau_3012_i1061(tree_3[21083:18072],tree_3[24095:21084],tree_3[27107:24096],tree_4[15059:12048],tree_4[18071:15060]);
csa_3012 csau_3012_i1062(tree_3[30119:27108],tree_3[33131:30120],tree_3[36143:33132],tree_4[21083:18072],tree_4[24095:21084]);
csa_3012 csau_3012_i1063(tree_3[39155:36144],tree_3[42167:39156],tree_3[45179:42168],tree_4[27107:24096],tree_4[30119:27108]);
csa_3012 csau_3012_i1064(tree_3[48191:45180],tree_3[51203:48192],tree_3[54215:51204],tree_4[33131:30120],tree_4[36143:33132]);
csa_3012 csau_3012_i1065(tree_3[57227:54216],tree_3[60239:57228],tree_3[63251:60240],tree_4[39155:36144],tree_4[42167:39156]);
csa_3012 csau_3012_i1066(tree_3[66263:63252],tree_3[69275:66264],tree_3[72287:69276],tree_4[45179:42168],tree_4[48191:45180]);
csa_3012 csau_3012_i1067(tree_3[75299:72288],tree_3[78311:75300],tree_3[81323:78312],tree_4[51203:48192],tree_4[54215:51204]);
csa_3012 csau_3012_i1068(tree_3[84335:81324],tree_3[87347:84336],tree_3[90359:87348],tree_4[57227:54216],tree_4[60239:57228]);
csa_3012 csau_3012_i1069(tree_3[93371:90360],tree_3[96383:93372],tree_3[99395:96384],tree_4[63251:60240],tree_4[66263:63252]);
csa_3012 csau_3012_i1070(tree_3[102407:99396],tree_3[105419:102408],tree_3[108431:105420],tree_4[69275:66264],tree_4[72287:69276]);
csa_3012 csau_3012_i1071(tree_3[111443:108432],tree_3[114455:111444],tree_3[117467:114456],tree_4[75299:72288],tree_4[78311:75300]);
csa_3012 csau_3012_i1072(tree_3[120479:117468],tree_3[123491:120480],tree_3[126503:123492],tree_4[81323:78312],tree_4[84335:81324]);
csa_3012 csau_3012_i1073(tree_3[129515:126504],tree_3[132527:129516],tree_3[135539:132528],tree_4[87347:84336],tree_4[90359:87348]);
csa_3012 csau_3012_i1074(tree_3[138551:135540],tree_3[141563:138552],tree_3[144575:141564],tree_4[93371:90360],tree_4[96383:93372]);
csa_3012 csau_3012_i1075(tree_3[147587:144576],tree_3[150599:147588],tree_3[153611:150600],tree_4[99395:96384],tree_4[102407:99396]);
csa_3012 csau_3012_i1076(tree_3[156623:153612],tree_3[159635:156624],tree_3[162647:159636],tree_4[105419:102408],tree_4[108431:105420]);
csa_3012 csau_3012_i1077(tree_3[165659:162648],tree_3[168671:165660],tree_3[171683:168672],tree_4[111443:108432],tree_4[114455:111444]);
csa_3012 csau_3012_i1078(tree_3[174695:171684],tree_3[177707:174696],tree_3[180719:177708],tree_4[117467:114456],tree_4[120479:117468]);
csa_3012 csau_3012_i1079(tree_3[183731:180720],tree_3[186743:183732],tree_3[189755:186744],tree_4[123491:120480],tree_4[126503:123492]);
csa_3012 csau_3012_i1080(tree_3[192767:189756],tree_3[195779:192768],tree_3[198791:195780],tree_4[129515:126504],tree_4[132527:129516]);
csa_3012 csau_3012_i1081(tree_3[201803:198792],tree_3[204815:201804],tree_3[207827:204816],tree_4[135539:132528],tree_4[138551:135540]);
csa_3012 csau_3012_i1082(tree_3[210839:207828],tree_3[213851:210840],tree_3[216863:213852],tree_4[141563:138552],tree_4[144575:141564]);
csa_3012 csau_3012_i1083(tree_3[219875:216864],tree_3[222887:219876],tree_3[225899:222888],tree_4[147587:144576],tree_4[150599:147588]);
csa_3012 csau_3012_i1084(tree_3[228911:225900],tree_3[231923:228912],tree_3[234935:231924],tree_4[153611:150600],tree_4[156623:153612]);
csa_3012 csau_3012_i1085(tree_3[237947:234936],tree_3[240959:237948],tree_3[243971:240960],tree_4[159635:156624],tree_4[162647:159636]);
csa_3012 csau_3012_i1086(tree_3[246983:243972],tree_3[249995:246984],tree_3[253007:249996],tree_4[165659:162648],tree_4[168671:165660]);
csa_3012 csau_3012_i1087(tree_3[256019:253008],tree_3[259031:256020],tree_3[262043:259032],tree_4[171683:168672],tree_4[174695:171684]);
csa_3012 csau_3012_i1088(tree_3[265055:262044],tree_3[268067:265056],tree_3[271079:268068],tree_4[177707:174696],tree_4[180719:177708]);
csa_3012 csau_3012_i1089(tree_3[274091:271080],tree_3[277103:274092],tree_3[280115:277104],tree_4[183731:180720],tree_4[186743:183732]);
csa_3012 csau_3012_i1090(tree_3[283127:280116],tree_3[286139:283128],tree_3[289151:286140],tree_4[189755:186744],tree_4[192767:189756]);
csa_3012 csau_3012_i1091(tree_3[292163:289152],tree_3[295175:292164],tree_3[298187:295176],tree_4[195779:192768],tree_4[198791:195780]);
csa_3012 csau_3012_i1092(tree_3[301199:298188],tree_3[304211:301200],tree_3[307223:304212],tree_4[201803:198792],tree_4[204815:201804]);
csa_3012 csau_3012_i1093(tree_3[310235:307224],tree_3[313247:310236],tree_3[316259:313248],tree_4[207827:204816],tree_4[210839:207828]);
csa_3012 csau_3012_i1094(tree_3[319271:316260],tree_3[322283:319272],tree_3[325295:322284],tree_4[213851:210840],tree_4[216863:213852]);
csa_3012 csau_3012_i1095(tree_3[328307:325296],tree_3[331319:328308],tree_3[334331:331320],tree_4[219875:216864],tree_4[222887:219876]);
csa_3012 csau_3012_i1096(tree_3[337343:334332],tree_3[340355:337344],tree_3[343367:340356],tree_4[225899:222888],tree_4[228911:225900]);
csa_3012 csau_3012_i1097(tree_3[346379:343368],tree_3[349391:346380],tree_3[352403:349392],tree_4[231923:228912],tree_4[234935:231924]);
csa_3012 csau_3012_i1098(tree_3[355415:352404],tree_3[358427:355416],tree_3[361439:358428],tree_4[237947:234936],tree_4[240959:237948]);
csa_3012 csau_3012_i1099(tree_3[364451:361440],tree_3[367463:364452],tree_3[370475:367464],tree_4[243971:240960],tree_4[246983:243972]);
csa_3012 csau_3012_i1100(tree_3[373487:370476],tree_3[376499:373488],tree_3[379511:376500],tree_4[249995:246984],tree_4[253007:249996]);
csa_3012 csau_3012_i1101(tree_3[382523:379512],tree_3[385535:382524],tree_3[388547:385536],tree_4[256019:253008],tree_4[259031:256020]);
csa_3012 csau_3012_i1102(tree_3[391559:388548],tree_3[394571:391560],tree_3[397583:394572],tree_4[262043:259032],tree_4[265055:262044]);
csa_3012 csau_3012_i1103(tree_3[400595:397584],tree_3[403607:400596],tree_3[406619:403608],tree_4[268067:265056],tree_4[271079:268068]);
csa_3012 csau_3012_i1104(tree_3[409631:406620],tree_3[412643:409632],tree_3[415655:412644],tree_4[274091:271080],tree_4[277103:274092]);
csa_3012 csau_3012_i1105(tree_3[418667:415656],tree_3[421679:418668],tree_3[424691:421680],tree_4[280115:277104],tree_4[283127:280116]);
csa_3012 csau_3012_i1106(tree_3[427703:424692],tree_3[430715:427704],tree_3[433727:430716],tree_4[286139:283128],tree_4[289151:286140]);
csa_3012 csau_3012_i1107(tree_3[436739:433728],tree_3[439751:436740],tree_3[442763:439752],tree_4[292163:289152],tree_4[295175:292164]);
csa_3012 csau_3012_i1108(tree_3[445775:442764],tree_3[448787:445776],tree_3[451799:448788],tree_4[298187:295176],tree_4[301199:298188]);
csa_3012 csau_3012_i1109(tree_3[454811:451800],tree_3[457823:454812],tree_3[460835:457824],tree_4[304211:301200],tree_4[307223:304212]);
csa_3012 csau_3012_i1110(tree_3[463847:460836],tree_3[466859:463848],tree_3[469871:466860],tree_4[310235:307224],tree_4[313247:310236]);
csa_3012 csau_3012_i1111(tree_3[472883:469872],tree_3[475895:472884],tree_3[478907:475896],tree_4[316259:313248],tree_4[319271:316260]);
csa_3012 csau_3012_i1112(tree_3[481919:478908],tree_3[484931:481920],tree_3[487943:484932],tree_4[322283:319272],tree_4[325295:322284]);
csa_3012 csau_3012_i1113(tree_3[490955:487944],tree_3[493967:490956],tree_3[496979:493968],tree_4[328307:325296],tree_4[331319:328308]);
csa_3012 csau_3012_i1114(tree_3[499991:496980],tree_3[503003:499992],tree_3[506015:503004],tree_4[334331:331320],tree_4[337343:334332]);
csa_3012 csau_3012_i1115(tree_3[509027:506016],tree_3[512039:509028],tree_3[515051:512040],tree_4[340355:337344],tree_4[343367:340356]);
csa_3012 csau_3012_i1116(tree_3[518063:515052],tree_3[521075:518064],tree_3[524087:521076],tree_4[346379:343368],tree_4[349391:346380]);
csa_3012 csau_3012_i1117(tree_3[527099:524088],tree_3[530111:527100],tree_3[533123:530112],tree_4[352403:349392],tree_4[355415:352404]);
csa_3012 csau_3012_i1118(tree_3[536135:533124],tree_3[539147:536136],tree_3[542159:539148],tree_4[358427:355416],tree_4[361439:358428]);
csa_3012 csau_3012_i1119(tree_3[545171:542160],tree_3[548183:545172],tree_3[551195:548184],tree_4[364451:361440],tree_4[367463:364452]);
csa_3012 csau_3012_i1120(tree_3[554207:551196],tree_3[557219:554208],tree_3[560231:557220],tree_4[370475:367464],tree_4[373487:370476]);
csa_3012 csau_3012_i1121(tree_3[563243:560232],tree_3[566255:563244],tree_3[569267:566256],tree_4[376499:373488],tree_4[379511:376500]);
csa_3012 csau_3012_i1122(tree_3[572279:569268],tree_3[575291:572280],tree_3[578303:575292],tree_4[382523:379512],tree_4[385535:382524]);
csa_3012 csau_3012_i1123(tree_3[581315:578304],tree_3[584327:581316],tree_3[587339:584328],tree_4[388547:385536],tree_4[391559:388548]);
csa_3012 csau_3012_i1124(tree_3[590351:587340],tree_3[593363:590352],tree_3[596375:593364],tree_4[394571:391560],tree_4[397583:394572]);
csa_3012 csau_3012_i1125(tree_3[599387:596376],tree_3[602399:599388],tree_3[605411:602400],tree_4[400595:397584],tree_4[403607:400596]);
csa_3012 csau_3012_i1126(tree_3[608423:605412],tree_3[611435:608424],tree_3[614447:611436],tree_4[406619:403608],tree_4[409631:406620]);
csa_3012 csau_3012_i1127(tree_3[617459:614448],tree_3[620471:617460],tree_3[623483:620472],tree_4[412643:409632],tree_4[415655:412644]);
csa_3012 csau_3012_i1128(tree_3[626495:623484],tree_3[629507:626496],tree_3[632519:629508],tree_4[418667:415656],tree_4[421679:418668]);
csa_3012 csau_3012_i1129(tree_3[635531:632520],tree_3[638543:635532],tree_3[641555:638544],tree_4[424691:421680],tree_4[427703:424692]);
csa_3012 csau_3012_i1130(tree_3[644567:641556],tree_3[647579:644568],tree_3[650591:647580],tree_4[430715:427704],tree_4[433727:430716]);
csa_3012 csau_3012_i1131(tree_3[653603:650592],tree_3[656615:653604],tree_3[659627:656616],tree_4[436739:433728],tree_4[439751:436740]);
csa_3012 csau_3012_i1132(tree_3[662639:659628],tree_3[665651:662640],tree_3[668663:665652],tree_4[442763:439752],tree_4[445775:442764]);
csa_3012 csau_3012_i1133(tree_3[671675:668664],tree_3[674687:671676],tree_3[677699:674688],tree_4[448787:445776],tree_4[451799:448788]);
csa_3012 csau_3012_i1134(tree_3[680711:677700],tree_3[683723:680712],tree_3[686735:683724],tree_4[454811:451800],tree_4[457823:454812]);
csa_3012 csau_3012_i1135(tree_3[689747:686736],tree_3[692759:689748],tree_3[695771:692760],tree_4[460835:457824],tree_4[463847:460836]);
csa_3012 csau_3012_i1136(tree_3[698783:695772],tree_3[701795:698784],tree_3[704807:701796],tree_4[466859:463848],tree_4[469871:466860]);
csa_3012 csau_3012_i1137(tree_3[707819:704808],tree_3[710831:707820],tree_3[713843:710832],tree_4[472883:469872],tree_4[475895:472884]);
csa_3012 csau_3012_i1138(tree_3[716855:713844],tree_3[719867:716856],tree_3[722879:719868],tree_4[478907:475896],tree_4[481919:478908]);
csa_3012 csau_3012_i1139(tree_3[725891:722880],tree_3[728903:725892],tree_3[731915:728904],tree_4[484931:481920],tree_4[487943:484932]);
csa_3012 csau_3012_i1140(tree_3[734927:731916],tree_3[737939:734928],tree_3[740951:737940],tree_4[490955:487944],tree_4[493967:490956]);
csa_3012 csau_3012_i1141(tree_3[743963:740952],tree_3[746975:743964],tree_3[749987:746976],tree_4[496979:493968],tree_4[499991:496980]);
csa_3012 csau_3012_i1142(tree_3[752999:749988],tree_3[756011:753000],tree_3[759023:756012],tree_4[503003:499992],tree_4[506015:503004]);
csa_3012 csau_3012_i1143(tree_3[762035:759024],tree_3[765047:762036],tree_3[768059:765048],tree_4[509027:506016],tree_4[512039:509028]);
csa_3012 csau_3012_i1144(tree_3[771071:768060],tree_3[774083:771072],tree_3[777095:774084],tree_4[515051:512040],tree_4[518063:515052]);
csa_3012 csau_3012_i1145(tree_3[780107:777096],tree_3[783119:780108],tree_3[786131:783120],tree_4[521075:518064],tree_4[524087:521076]);
csa_3012 csau_3012_i1146(tree_3[789143:786132],tree_3[792155:789144],tree_3[795167:792156],tree_4[527099:524088],tree_4[530111:527100]);
csa_3012 csau_3012_i1147(tree_3[798179:795168],tree_3[801191:798180],tree_3[804203:801192],tree_4[533123:530112],tree_4[536135:533124]);
csa_3012 csau_3012_i1148(tree_3[807215:804204],tree_3[810227:807216],tree_3[813239:810228],tree_4[539147:536136],tree_4[542159:539148]);
csa_3012 csau_3012_i1149(tree_3[816251:813240],tree_3[819263:816252],tree_3[822275:819264],tree_4[545171:542160],tree_4[548183:545172]);
csa_3012 csau_3012_i1150(tree_3[825287:822276],tree_3[828299:825288],tree_3[831311:828300],tree_4[551195:548184],tree_4[554207:551196]);
csa_3012 csau_3012_i1151(tree_3[834323:831312],tree_3[837335:834324],tree_3[840347:837336],tree_4[557219:554208],tree_4[560231:557220]);
csa_3012 csau_3012_i1152(tree_3[843359:840348],tree_3[846371:843360],tree_3[849383:846372],tree_4[563243:560232],tree_4[566255:563244]);
csa_3012 csau_3012_i1153(tree_3[852395:849384],tree_3[855407:852396],tree_3[858419:855408],tree_4[569267:566256],tree_4[572279:569268]);
csa_3012 csau_3012_i1154(tree_3[861431:858420],tree_3[864443:861432],tree_3[867455:864444],tree_4[575291:572280],tree_4[578303:575292]);
csa_3012 csau_3012_i1155(tree_3[870467:867456],tree_3[873479:870468],tree_3[876491:873480],tree_4[581315:578304],tree_4[584327:581316]);
csa_3012 csau_3012_i1156(tree_3[879503:876492],tree_3[882515:879504],tree_3[885527:882516],tree_4[587339:584328],tree_4[590351:587340]);
csa_3012 csau_3012_i1157(tree_3[888539:885528],tree_3[891551:888540],tree_3[894563:891552],tree_4[593363:590352],tree_4[596375:593364]);
csa_3012 csau_3012_i1158(tree_3[897575:894564],tree_3[900587:897576],tree_3[903599:900588],tree_4[599387:596376],tree_4[602399:599388]);
csa_3012 csau_3012_i1159(tree_3[906611:903600],tree_3[909623:906612],tree_3[912635:909624],tree_4[605411:602400],tree_4[608423:605412]);
csa_3012 csau_3012_i1160(tree_3[915647:912636],tree_3[918659:915648],tree_3[921671:918660],tree_4[611435:608424],tree_4[614447:611436]);
csa_3012 csau_3012_i1161(tree_3[924683:921672],tree_3[927695:924684],tree_3[930707:927696],tree_4[617459:614448],tree_4[620471:617460]);
csa_3012 csau_3012_i1162(tree_3[933719:930708],tree_3[936731:933720],tree_3[939743:936732],tree_4[623483:620472],tree_4[626495:623484]);
csa_3012 csau_3012_i1163(tree_3[942755:939744],tree_3[945767:942756],tree_3[948779:945768],tree_4[629507:626496],tree_4[632519:629508]);
csa_3012 csau_3012_i1164(tree_3[951791:948780],tree_3[954803:951792],tree_3[957815:954804],tree_4[635531:632520],tree_4[638543:635532]);
csa_3012 csau_3012_i1165(tree_3[960827:957816],tree_3[963839:960828],tree_3[966851:963840],tree_4[641555:638544],tree_4[644567:641556]);
csa_3012 csau_3012_i1166(tree_3[969863:966852],tree_3[972875:969864],tree_3[975887:972876],tree_4[647579:644568],tree_4[650591:647580]);
csa_3012 csau_3012_i1167(tree_3[978899:975888],tree_3[981911:978900],tree_3[984923:981912],tree_4[653603:650592],tree_4[656615:653604]);
csa_3012 csau_3012_i1168(tree_3[987935:984924],tree_3[990947:987936],tree_3[993959:990948],tree_4[659627:656616],tree_4[662639:659628]);
csa_3012 csau_3012_i1169(tree_3[996971:993960],tree_3[999983:996972],tree_3[1002995:999984],tree_4[665651:662640],tree_4[668663:665652]);
csa_3012 csau_3012_i1170(tree_3[1006007:1002996],tree_3[1009019:1006008],tree_3[1012031:1009020],tree_4[671675:668664],tree_4[674687:671676]);
csa_3012 csau_3012_i1171(tree_3[1015043:1012032],tree_3[1018055:1015044],tree_3[1021067:1018056],tree_4[677699:674688],tree_4[680711:677700]);
csa_3012 csau_3012_i1172(tree_3[1024079:1021068],tree_3[1027091:1024080],tree_3[1030103:1027092],tree_4[683723:680712],tree_4[686735:683724]);
csa_3012 csau_3012_i1173(tree_3[1033115:1030104],tree_3[1036127:1033116],tree_3[1039139:1036128],tree_4[689747:686736],tree_4[692759:689748]);
csa_3012 csau_3012_i1174(tree_3[1042151:1039140],tree_3[1045163:1042152],tree_3[1048175:1045164],tree_4[695771:692760],tree_4[698783:695772]);
csa_3012 csau_3012_i1175(tree_3[1051187:1048176],tree_3[1054199:1051188],tree_3[1057211:1054200],tree_4[701795:698784],tree_4[704807:701796]);
csa_3012 csau_3012_i1176(tree_3[1060223:1057212],tree_3[1063235:1060224],tree_3[1066247:1063236],tree_4[707819:704808],tree_4[710831:707820]);
csa_3012 csau_3012_i1177(tree_3[1069259:1066248],tree_3[1072271:1069260],tree_3[1075283:1072272],tree_4[713843:710832],tree_4[716855:713844]);
csa_3012 csau_3012_i1178(tree_3[1078295:1075284],tree_3[1081307:1078296],tree_3[1084319:1081308],tree_4[719867:716856],tree_4[722879:719868]);
csa_3012 csau_3012_i1179(tree_3[1087331:1084320],tree_3[1090343:1087332],tree_3[1093355:1090344],tree_4[725891:722880],tree_4[728903:725892]);
csa_3012 csau_3012_i1180(tree_3[1096367:1093356],tree_3[1099379:1096368],tree_3[1102391:1099380],tree_4[731915:728904],tree_4[734927:731916]);
csa_3012 csau_3012_i1181(tree_3[1105403:1102392],tree_3[1108415:1105404],tree_3[1111427:1108416],tree_4[737939:734928],tree_4[740951:737940]);
csa_3012 csau_3012_i1182(tree_3[1114439:1111428],tree_3[1117451:1114440],tree_3[1120463:1117452],tree_4[743963:740952],tree_4[746975:743964]);
csa_3012 csau_3012_i1183(tree_3[1123475:1120464],tree_3[1126487:1123476],tree_3[1129499:1126488],tree_4[749987:746976],tree_4[752999:749988]);
csa_3012 csau_3012_i1184(tree_3[1132511:1129500],tree_3[1135523:1132512],tree_3[1138535:1135524],tree_4[756011:753000],tree_4[759023:756012]);
csa_3012 csau_3012_i1185(tree_3[1141547:1138536],tree_3[1144559:1141548],tree_3[1147571:1144560],tree_4[762035:759024],tree_4[765047:762036]);
csa_3012 csau_3012_i1186(tree_3[1150583:1147572],tree_3[1153595:1150584],tree_3[1156607:1153596],tree_4[768059:765048],tree_4[771071:768060]);
csa_3012 csau_3012_i1187(tree_3[1159619:1156608],tree_3[1162631:1159620],tree_3[1165643:1162632],tree_4[774083:771072],tree_4[777095:774084]);
csa_3012 csau_3012_i1188(tree_3[1168655:1165644],tree_3[1171667:1168656],tree_3[1174679:1171668],tree_4[780107:777096],tree_4[783119:780108]);
csa_3012 csau_3012_i1189(tree_3[1177691:1174680],tree_3[1180703:1177692],tree_3[1183715:1180704],tree_4[786131:783120],tree_4[789143:786132]);
csa_3012 csau_3012_i1190(tree_3[1186727:1183716],tree_3[1189739:1186728],tree_3[1192751:1189740],tree_4[792155:789144],tree_4[795167:792156]);
csa_3012 csau_3012_i1191(tree_3[1195763:1192752],tree_3[1198775:1195764],tree_3[1201787:1198776],tree_4[798179:795168],tree_4[801191:798180]);
csa_3012 csau_3012_i1192(tree_3[1204799:1201788],tree_3[1207811:1204800],tree_3[1210823:1207812],tree_4[804203:801192],tree_4[807215:804204]);
csa_3012 csau_3012_i1193(tree_3[1213835:1210824],tree_3[1216847:1213836],tree_3[1219859:1216848],tree_4[810227:807216],tree_4[813239:810228]);
csa_3012 csau_3012_i1194(tree_3[1222871:1219860],tree_3[1225883:1222872],tree_3[1228895:1225884],tree_4[816251:813240],tree_4[819263:816252]);
csa_3012 csau_3012_i1195(tree_3[1231907:1228896],tree_3[1234919:1231908],tree_3[1237931:1234920],tree_4[822275:819264],tree_4[825287:822276]);
csa_3012 csau_3012_i1196(tree_3[1240943:1237932],tree_3[1243955:1240944],tree_3[1246967:1243956],tree_4[828299:825288],tree_4[831311:828300]);
csa_3012 csau_3012_i1197(tree_3[1249979:1246968],tree_3[1252991:1249980],tree_3[1256003:1252992],tree_4[834323:831312],tree_4[837335:834324]);
csa_3012 csau_3012_i1198(tree_3[1259015:1256004],tree_3[1262027:1259016],tree_3[1265039:1262028],tree_4[840347:837336],tree_4[843359:840348]);
csa_3012 csau_3012_i1199(tree_3[1268051:1265040],tree_3[1271063:1268052],tree_3[1274075:1271064],tree_4[846371:843360],tree_4[849383:846372]);
csa_3012 csau_3012_i1200(tree_3[1277087:1274076],tree_3[1280099:1277088],tree_3[1283111:1280100],tree_4[852395:849384],tree_4[855407:852396]);
csa_3012 csau_3012_i1201(tree_3[1286123:1283112],tree_3[1289135:1286124],tree_3[1292147:1289136],tree_4[858419:855408],tree_4[861431:858420]);
csa_3012 csau_3012_i1202(tree_3[1295159:1292148],tree_3[1298171:1295160],tree_3[1301183:1298172],tree_4[864443:861432],tree_4[867455:864444]);
csa_3012 csau_3012_i1203(tree_3[1304195:1301184],tree_3[1307207:1304196],tree_3[1310219:1307208],tree_4[870467:867456],tree_4[873479:870468]);
csa_3012 csau_3012_i1204(tree_3[1313231:1310220],tree_3[1316243:1313232],tree_3[1319255:1316244],tree_4[876491:873480],tree_4[879503:876492]);
csa_3012 csau_3012_i1205(tree_3[1322267:1319256],tree_3[1325279:1322268],tree_3[1328291:1325280],tree_4[882515:879504],tree_4[885527:882516]);
csa_3012 csau_3012_i1206(tree_3[1331303:1328292],tree_3[1334315:1331304],tree_3[1337327:1334316],tree_4[888539:885528],tree_4[891551:888540]);
csa_3012 csau_3012_i1207(tree_3[1340339:1337328],tree_3[1343351:1340340],tree_3[1346363:1343352],tree_4[894563:891552],tree_4[897575:894564]);
// layer-5
csa_3012 csau_3012_i1208(tree_4[3011:0],tree_4[6023:3012],tree_4[9035:6024],tree_5[3011:0],tree_5[6023:3012]);
csa_3012 csau_3012_i1209(tree_4[12047:9036],tree_4[15059:12048],tree_4[18071:15060],tree_5[9035:6024],tree_5[12047:9036]);
csa_3012 csau_3012_i1210(tree_4[21083:18072],tree_4[24095:21084],tree_4[27107:24096],tree_5[15059:12048],tree_5[18071:15060]);
csa_3012 csau_3012_i1211(tree_4[30119:27108],tree_4[33131:30120],tree_4[36143:33132],tree_5[21083:18072],tree_5[24095:21084]);
csa_3012 csau_3012_i1212(tree_4[39155:36144],tree_4[42167:39156],tree_4[45179:42168],tree_5[27107:24096],tree_5[30119:27108]);
csa_3012 csau_3012_i1213(tree_4[48191:45180],tree_4[51203:48192],tree_4[54215:51204],tree_5[33131:30120],tree_5[36143:33132]);
csa_3012 csau_3012_i1214(tree_4[57227:54216],tree_4[60239:57228],tree_4[63251:60240],tree_5[39155:36144],tree_5[42167:39156]);
csa_3012 csau_3012_i1215(tree_4[66263:63252],tree_4[69275:66264],tree_4[72287:69276],tree_5[45179:42168],tree_5[48191:45180]);
csa_3012 csau_3012_i1216(tree_4[75299:72288],tree_4[78311:75300],tree_4[81323:78312],tree_5[51203:48192],tree_5[54215:51204]);
csa_3012 csau_3012_i1217(tree_4[84335:81324],tree_4[87347:84336],tree_4[90359:87348],tree_5[57227:54216],tree_5[60239:57228]);
csa_3012 csau_3012_i1218(tree_4[93371:90360],tree_4[96383:93372],tree_4[99395:96384],tree_5[63251:60240],tree_5[66263:63252]);
csa_3012 csau_3012_i1219(tree_4[102407:99396],tree_4[105419:102408],tree_4[108431:105420],tree_5[69275:66264],tree_5[72287:69276]);
csa_3012 csau_3012_i1220(tree_4[111443:108432],tree_4[114455:111444],tree_4[117467:114456],tree_5[75299:72288],tree_5[78311:75300]);
csa_3012 csau_3012_i1221(tree_4[120479:117468],tree_4[123491:120480],tree_4[126503:123492],tree_5[81323:78312],tree_5[84335:81324]);
csa_3012 csau_3012_i1222(tree_4[129515:126504],tree_4[132527:129516],tree_4[135539:132528],tree_5[87347:84336],tree_5[90359:87348]);
csa_3012 csau_3012_i1223(tree_4[138551:135540],tree_4[141563:138552],tree_4[144575:141564],tree_5[93371:90360],tree_5[96383:93372]);
csa_3012 csau_3012_i1224(tree_4[147587:144576],tree_4[150599:147588],tree_4[153611:150600],tree_5[99395:96384],tree_5[102407:99396]);
csa_3012 csau_3012_i1225(tree_4[156623:153612],tree_4[159635:156624],tree_4[162647:159636],tree_5[105419:102408],tree_5[108431:105420]);
csa_3012 csau_3012_i1226(tree_4[165659:162648],tree_4[168671:165660],tree_4[171683:168672],tree_5[111443:108432],tree_5[114455:111444]);
csa_3012 csau_3012_i1227(tree_4[174695:171684],tree_4[177707:174696],tree_4[180719:177708],tree_5[117467:114456],tree_5[120479:117468]);
csa_3012 csau_3012_i1228(tree_4[183731:180720],tree_4[186743:183732],tree_4[189755:186744],tree_5[123491:120480],tree_5[126503:123492]);
csa_3012 csau_3012_i1229(tree_4[192767:189756],tree_4[195779:192768],tree_4[198791:195780],tree_5[129515:126504],tree_5[132527:129516]);
csa_3012 csau_3012_i1230(tree_4[201803:198792],tree_4[204815:201804],tree_4[207827:204816],tree_5[135539:132528],tree_5[138551:135540]);
csa_3012 csau_3012_i1231(tree_4[210839:207828],tree_4[213851:210840],tree_4[216863:213852],tree_5[141563:138552],tree_5[144575:141564]);
csa_3012 csau_3012_i1232(tree_4[219875:216864],tree_4[222887:219876],tree_4[225899:222888],tree_5[147587:144576],tree_5[150599:147588]);
csa_3012 csau_3012_i1233(tree_4[228911:225900],tree_4[231923:228912],tree_4[234935:231924],tree_5[153611:150600],tree_5[156623:153612]);
csa_3012 csau_3012_i1234(tree_4[237947:234936],tree_4[240959:237948],tree_4[243971:240960],tree_5[159635:156624],tree_5[162647:159636]);
csa_3012 csau_3012_i1235(tree_4[246983:243972],tree_4[249995:246984],tree_4[253007:249996],tree_5[165659:162648],tree_5[168671:165660]);
csa_3012 csau_3012_i1236(tree_4[256019:253008],tree_4[259031:256020],tree_4[262043:259032],tree_5[171683:168672],tree_5[174695:171684]);
csa_3012 csau_3012_i1237(tree_4[265055:262044],tree_4[268067:265056],tree_4[271079:268068],tree_5[177707:174696],tree_5[180719:177708]);
csa_3012 csau_3012_i1238(tree_4[274091:271080],tree_4[277103:274092],tree_4[280115:277104],tree_5[183731:180720],tree_5[186743:183732]);
csa_3012 csau_3012_i1239(tree_4[283127:280116],tree_4[286139:283128],tree_4[289151:286140],tree_5[189755:186744],tree_5[192767:189756]);
csa_3012 csau_3012_i1240(tree_4[292163:289152],tree_4[295175:292164],tree_4[298187:295176],tree_5[195779:192768],tree_5[198791:195780]);
csa_3012 csau_3012_i1241(tree_4[301199:298188],tree_4[304211:301200],tree_4[307223:304212],tree_5[201803:198792],tree_5[204815:201804]);
csa_3012 csau_3012_i1242(tree_4[310235:307224],tree_4[313247:310236],tree_4[316259:313248],tree_5[207827:204816],tree_5[210839:207828]);
csa_3012 csau_3012_i1243(tree_4[319271:316260],tree_4[322283:319272],tree_4[325295:322284],tree_5[213851:210840],tree_5[216863:213852]);
csa_3012 csau_3012_i1244(tree_4[328307:325296],tree_4[331319:328308],tree_4[334331:331320],tree_5[219875:216864],tree_5[222887:219876]);
csa_3012 csau_3012_i1245(tree_4[337343:334332],tree_4[340355:337344],tree_4[343367:340356],tree_5[225899:222888],tree_5[228911:225900]);
csa_3012 csau_3012_i1246(tree_4[346379:343368],tree_4[349391:346380],tree_4[352403:349392],tree_5[231923:228912],tree_5[234935:231924]);
csa_3012 csau_3012_i1247(tree_4[355415:352404],tree_4[358427:355416],tree_4[361439:358428],tree_5[237947:234936],tree_5[240959:237948]);
csa_3012 csau_3012_i1248(tree_4[364451:361440],tree_4[367463:364452],tree_4[370475:367464],tree_5[243971:240960],tree_5[246983:243972]);
csa_3012 csau_3012_i1249(tree_4[373487:370476],tree_4[376499:373488],tree_4[379511:376500],tree_5[249995:246984],tree_5[253007:249996]);
csa_3012 csau_3012_i1250(tree_4[382523:379512],tree_4[385535:382524],tree_4[388547:385536],tree_5[256019:253008],tree_5[259031:256020]);
csa_3012 csau_3012_i1251(tree_4[391559:388548],tree_4[394571:391560],tree_4[397583:394572],tree_5[262043:259032],tree_5[265055:262044]);
csa_3012 csau_3012_i1252(tree_4[400595:397584],tree_4[403607:400596],tree_4[406619:403608],tree_5[268067:265056],tree_5[271079:268068]);
csa_3012 csau_3012_i1253(tree_4[409631:406620],tree_4[412643:409632],tree_4[415655:412644],tree_5[274091:271080],tree_5[277103:274092]);
csa_3012 csau_3012_i1254(tree_4[418667:415656],tree_4[421679:418668],tree_4[424691:421680],tree_5[280115:277104],tree_5[283127:280116]);
csa_3012 csau_3012_i1255(tree_4[427703:424692],tree_4[430715:427704],tree_4[433727:430716],tree_5[286139:283128],tree_5[289151:286140]);
csa_3012 csau_3012_i1256(tree_4[436739:433728],tree_4[439751:436740],tree_4[442763:439752],tree_5[292163:289152],tree_5[295175:292164]);
csa_3012 csau_3012_i1257(tree_4[445775:442764],tree_4[448787:445776],tree_4[451799:448788],tree_5[298187:295176],tree_5[301199:298188]);
csa_3012 csau_3012_i1258(tree_4[454811:451800],tree_4[457823:454812],tree_4[460835:457824],tree_5[304211:301200],tree_5[307223:304212]);
csa_3012 csau_3012_i1259(tree_4[463847:460836],tree_4[466859:463848],tree_4[469871:466860],tree_5[310235:307224],tree_5[313247:310236]);
csa_3012 csau_3012_i1260(tree_4[472883:469872],tree_4[475895:472884],tree_4[478907:475896],tree_5[316259:313248],tree_5[319271:316260]);
csa_3012 csau_3012_i1261(tree_4[481919:478908],tree_4[484931:481920],tree_4[487943:484932],tree_5[322283:319272],tree_5[325295:322284]);
csa_3012 csau_3012_i1262(tree_4[490955:487944],tree_4[493967:490956],tree_4[496979:493968],tree_5[328307:325296],tree_5[331319:328308]);
csa_3012 csau_3012_i1263(tree_4[499991:496980],tree_4[503003:499992],tree_4[506015:503004],tree_5[334331:331320],tree_5[337343:334332]);
csa_3012 csau_3012_i1264(tree_4[509027:506016],tree_4[512039:509028],tree_4[515051:512040],tree_5[340355:337344],tree_5[343367:340356]);
csa_3012 csau_3012_i1265(tree_4[518063:515052],tree_4[521075:518064],tree_4[524087:521076],tree_5[346379:343368],tree_5[349391:346380]);
csa_3012 csau_3012_i1266(tree_4[527099:524088],tree_4[530111:527100],tree_4[533123:530112],tree_5[352403:349392],tree_5[355415:352404]);
csa_3012 csau_3012_i1267(tree_4[536135:533124],tree_4[539147:536136],tree_4[542159:539148],tree_5[358427:355416],tree_5[361439:358428]);
csa_3012 csau_3012_i1268(tree_4[545171:542160],tree_4[548183:545172],tree_4[551195:548184],tree_5[364451:361440],tree_5[367463:364452]);
csa_3012 csau_3012_i1269(tree_4[554207:551196],tree_4[557219:554208],tree_4[560231:557220],tree_5[370475:367464],tree_5[373487:370476]);
csa_3012 csau_3012_i1270(tree_4[563243:560232],tree_4[566255:563244],tree_4[569267:566256],tree_5[376499:373488],tree_5[379511:376500]);
csa_3012 csau_3012_i1271(tree_4[572279:569268],tree_4[575291:572280],tree_4[578303:575292],tree_5[382523:379512],tree_5[385535:382524]);
csa_3012 csau_3012_i1272(tree_4[581315:578304],tree_4[584327:581316],tree_4[587339:584328],tree_5[388547:385536],tree_5[391559:388548]);
csa_3012 csau_3012_i1273(tree_4[590351:587340],tree_4[593363:590352],tree_4[596375:593364],tree_5[394571:391560],tree_5[397583:394572]);
csa_3012 csau_3012_i1274(tree_4[599387:596376],tree_4[602399:599388],tree_4[605411:602400],tree_5[400595:397584],tree_5[403607:400596]);
csa_3012 csau_3012_i1275(tree_4[608423:605412],tree_4[611435:608424],tree_4[614447:611436],tree_5[406619:403608],tree_5[409631:406620]);
csa_3012 csau_3012_i1276(tree_4[617459:614448],tree_4[620471:617460],tree_4[623483:620472],tree_5[412643:409632],tree_5[415655:412644]);
csa_3012 csau_3012_i1277(tree_4[626495:623484],tree_4[629507:626496],tree_4[632519:629508],tree_5[418667:415656],tree_5[421679:418668]);
csa_3012 csau_3012_i1278(tree_4[635531:632520],tree_4[638543:635532],tree_4[641555:638544],tree_5[424691:421680],tree_5[427703:424692]);
csa_3012 csau_3012_i1279(tree_4[644567:641556],tree_4[647579:644568],tree_4[650591:647580],tree_5[430715:427704],tree_5[433727:430716]);
csa_3012 csau_3012_i1280(tree_4[653603:650592],tree_4[656615:653604],tree_4[659627:656616],tree_5[436739:433728],tree_5[439751:436740]);
csa_3012 csau_3012_i1281(tree_4[662639:659628],tree_4[665651:662640],tree_4[668663:665652],tree_5[442763:439752],tree_5[445775:442764]);
csa_3012 csau_3012_i1282(tree_4[671675:668664],tree_4[674687:671676],tree_4[677699:674688],tree_5[448787:445776],tree_5[451799:448788]);
csa_3012 csau_3012_i1283(tree_4[680711:677700],tree_4[683723:680712],tree_4[686735:683724],tree_5[454811:451800],tree_5[457823:454812]);
csa_3012 csau_3012_i1284(tree_4[689747:686736],tree_4[692759:689748],tree_4[695771:692760],tree_5[460835:457824],tree_5[463847:460836]);
csa_3012 csau_3012_i1285(tree_4[698783:695772],tree_4[701795:698784],tree_4[704807:701796],tree_5[466859:463848],tree_5[469871:466860]);
csa_3012 csau_3012_i1286(tree_4[707819:704808],tree_4[710831:707820],tree_4[713843:710832],tree_5[472883:469872],tree_5[475895:472884]);
csa_3012 csau_3012_i1287(tree_4[716855:713844],tree_4[719867:716856],tree_4[722879:719868],tree_5[478907:475896],tree_5[481919:478908]);
csa_3012 csau_3012_i1288(tree_4[725891:722880],tree_4[728903:725892],tree_4[731915:728904],tree_5[484931:481920],tree_5[487943:484932]);
csa_3012 csau_3012_i1289(tree_4[734927:731916],tree_4[737939:734928],tree_4[740951:737940],tree_5[490955:487944],tree_5[493967:490956]);
csa_3012 csau_3012_i1290(tree_4[743963:740952],tree_4[746975:743964],tree_4[749987:746976],tree_5[496979:493968],tree_5[499991:496980]);
csa_3012 csau_3012_i1291(tree_4[752999:749988],tree_4[756011:753000],tree_4[759023:756012],tree_5[503003:499992],tree_5[506015:503004]);
csa_3012 csau_3012_i1292(tree_4[762035:759024],tree_4[765047:762036],tree_4[768059:765048],tree_5[509027:506016],tree_5[512039:509028]);
csa_3012 csau_3012_i1293(tree_4[771071:768060],tree_4[774083:771072],tree_4[777095:774084],tree_5[515051:512040],tree_5[518063:515052]);
csa_3012 csau_3012_i1294(tree_4[780107:777096],tree_4[783119:780108],tree_4[786131:783120],tree_5[521075:518064],tree_5[524087:521076]);
csa_3012 csau_3012_i1295(tree_4[789143:786132],tree_4[792155:789144],tree_4[795167:792156],tree_5[527099:524088],tree_5[530111:527100]);
csa_3012 csau_3012_i1296(tree_4[798179:795168],tree_4[801191:798180],tree_4[804203:801192],tree_5[533123:530112],tree_5[536135:533124]);
csa_3012 csau_3012_i1297(tree_4[807215:804204],tree_4[810227:807216],tree_4[813239:810228],tree_5[539147:536136],tree_5[542159:539148]);
csa_3012 csau_3012_i1298(tree_4[816251:813240],tree_4[819263:816252],tree_4[822275:819264],tree_5[545171:542160],tree_5[548183:545172]);
csa_3012 csau_3012_i1299(tree_4[825287:822276],tree_4[828299:825288],tree_4[831311:828300],tree_5[551195:548184],tree_5[554207:551196]);
csa_3012 csau_3012_i1300(tree_4[834323:831312],tree_4[837335:834324],tree_4[840347:837336],tree_5[557219:554208],tree_5[560231:557220]);
csa_3012 csau_3012_i1301(tree_4[843359:840348],tree_4[846371:843360],tree_4[849383:846372],tree_5[563243:560232],tree_5[566255:563244]);
csa_3012 csau_3012_i1302(tree_4[852395:849384],tree_4[855407:852396],tree_4[858419:855408],tree_5[569267:566256],tree_5[572279:569268]);
csa_3012 csau_3012_i1303(tree_4[861431:858420],tree_4[864443:861432],tree_4[867455:864444],tree_5[575291:572280],tree_5[578303:575292]);
csa_3012 csau_3012_i1304(tree_4[870467:867456],tree_4[873479:870468],tree_4[876491:873480],tree_5[581315:578304],tree_5[584327:581316]);
csa_3012 csau_3012_i1305(tree_4[879503:876492],tree_4[882515:879504],tree_4[885527:882516],tree_5[587339:584328],tree_5[590351:587340]);
csa_3012 csau_3012_i1306(tree_4[888539:885528],tree_4[891551:888540],tree_4[894563:891552],tree_5[593363:590352],tree_5[596375:593364]);
assign tree_5[599387:596376] = tree_4[897575:894564];
// layer-6
csa_3012 csau_3012_i1307(tree_5[3011:0],tree_5[6023:3012],tree_5[9035:6024],tree_6[3011:0],tree_6[6023:3012]);
csa_3012 csau_3012_i1308(tree_5[12047:9036],tree_5[15059:12048],tree_5[18071:15060],tree_6[9035:6024],tree_6[12047:9036]);
csa_3012 csau_3012_i1309(tree_5[21083:18072],tree_5[24095:21084],tree_5[27107:24096],tree_6[15059:12048],tree_6[18071:15060]);
csa_3012 csau_3012_i1310(tree_5[30119:27108],tree_5[33131:30120],tree_5[36143:33132],tree_6[21083:18072],tree_6[24095:21084]);
csa_3012 csau_3012_i1311(tree_5[39155:36144],tree_5[42167:39156],tree_5[45179:42168],tree_6[27107:24096],tree_6[30119:27108]);
csa_3012 csau_3012_i1312(tree_5[48191:45180],tree_5[51203:48192],tree_5[54215:51204],tree_6[33131:30120],tree_6[36143:33132]);
csa_3012 csau_3012_i1313(tree_5[57227:54216],tree_5[60239:57228],tree_5[63251:60240],tree_6[39155:36144],tree_6[42167:39156]);
csa_3012 csau_3012_i1314(tree_5[66263:63252],tree_5[69275:66264],tree_5[72287:69276],tree_6[45179:42168],tree_6[48191:45180]);
csa_3012 csau_3012_i1315(tree_5[75299:72288],tree_5[78311:75300],tree_5[81323:78312],tree_6[51203:48192],tree_6[54215:51204]);
csa_3012 csau_3012_i1316(tree_5[84335:81324],tree_5[87347:84336],tree_5[90359:87348],tree_6[57227:54216],tree_6[60239:57228]);
csa_3012 csau_3012_i1317(tree_5[93371:90360],tree_5[96383:93372],tree_5[99395:96384],tree_6[63251:60240],tree_6[66263:63252]);
csa_3012 csau_3012_i1318(tree_5[102407:99396],tree_5[105419:102408],tree_5[108431:105420],tree_6[69275:66264],tree_6[72287:69276]);
csa_3012 csau_3012_i1319(tree_5[111443:108432],tree_5[114455:111444],tree_5[117467:114456],tree_6[75299:72288],tree_6[78311:75300]);
csa_3012 csau_3012_i1320(tree_5[120479:117468],tree_5[123491:120480],tree_5[126503:123492],tree_6[81323:78312],tree_6[84335:81324]);
csa_3012 csau_3012_i1321(tree_5[129515:126504],tree_5[132527:129516],tree_5[135539:132528],tree_6[87347:84336],tree_6[90359:87348]);
csa_3012 csau_3012_i1322(tree_5[138551:135540],tree_5[141563:138552],tree_5[144575:141564],tree_6[93371:90360],tree_6[96383:93372]);
csa_3012 csau_3012_i1323(tree_5[147587:144576],tree_5[150599:147588],tree_5[153611:150600],tree_6[99395:96384],tree_6[102407:99396]);
csa_3012 csau_3012_i1324(tree_5[156623:153612],tree_5[159635:156624],tree_5[162647:159636],tree_6[105419:102408],tree_6[108431:105420]);
csa_3012 csau_3012_i1325(tree_5[165659:162648],tree_5[168671:165660],tree_5[171683:168672],tree_6[111443:108432],tree_6[114455:111444]);
csa_3012 csau_3012_i1326(tree_5[174695:171684],tree_5[177707:174696],tree_5[180719:177708],tree_6[117467:114456],tree_6[120479:117468]);
csa_3012 csau_3012_i1327(tree_5[183731:180720],tree_5[186743:183732],tree_5[189755:186744],tree_6[123491:120480],tree_6[126503:123492]);
csa_3012 csau_3012_i1328(tree_5[192767:189756],tree_5[195779:192768],tree_5[198791:195780],tree_6[129515:126504],tree_6[132527:129516]);
csa_3012 csau_3012_i1329(tree_5[201803:198792],tree_5[204815:201804],tree_5[207827:204816],tree_6[135539:132528],tree_6[138551:135540]);
csa_3012 csau_3012_i1330(tree_5[210839:207828],tree_5[213851:210840],tree_5[216863:213852],tree_6[141563:138552],tree_6[144575:141564]);
csa_3012 csau_3012_i1331(tree_5[219875:216864],tree_5[222887:219876],tree_5[225899:222888],tree_6[147587:144576],tree_6[150599:147588]);
csa_3012 csau_3012_i1332(tree_5[228911:225900],tree_5[231923:228912],tree_5[234935:231924],tree_6[153611:150600],tree_6[156623:153612]);
csa_3012 csau_3012_i1333(tree_5[237947:234936],tree_5[240959:237948],tree_5[243971:240960],tree_6[159635:156624],tree_6[162647:159636]);
csa_3012 csau_3012_i1334(tree_5[246983:243972],tree_5[249995:246984],tree_5[253007:249996],tree_6[165659:162648],tree_6[168671:165660]);
csa_3012 csau_3012_i1335(tree_5[256019:253008],tree_5[259031:256020],tree_5[262043:259032],tree_6[171683:168672],tree_6[174695:171684]);
csa_3012 csau_3012_i1336(tree_5[265055:262044],tree_5[268067:265056],tree_5[271079:268068],tree_6[177707:174696],tree_6[180719:177708]);
csa_3012 csau_3012_i1337(tree_5[274091:271080],tree_5[277103:274092],tree_5[280115:277104],tree_6[183731:180720],tree_6[186743:183732]);
csa_3012 csau_3012_i1338(tree_5[283127:280116],tree_5[286139:283128],tree_5[289151:286140],tree_6[189755:186744],tree_6[192767:189756]);
csa_3012 csau_3012_i1339(tree_5[292163:289152],tree_5[295175:292164],tree_5[298187:295176],tree_6[195779:192768],tree_6[198791:195780]);
csa_3012 csau_3012_i1340(tree_5[301199:298188],tree_5[304211:301200],tree_5[307223:304212],tree_6[201803:198792],tree_6[204815:201804]);
csa_3012 csau_3012_i1341(tree_5[310235:307224],tree_5[313247:310236],tree_5[316259:313248],tree_6[207827:204816],tree_6[210839:207828]);
csa_3012 csau_3012_i1342(tree_5[319271:316260],tree_5[322283:319272],tree_5[325295:322284],tree_6[213851:210840],tree_6[216863:213852]);
csa_3012 csau_3012_i1343(tree_5[328307:325296],tree_5[331319:328308],tree_5[334331:331320],tree_6[219875:216864],tree_6[222887:219876]);
csa_3012 csau_3012_i1344(tree_5[337343:334332],tree_5[340355:337344],tree_5[343367:340356],tree_6[225899:222888],tree_6[228911:225900]);
csa_3012 csau_3012_i1345(tree_5[346379:343368],tree_5[349391:346380],tree_5[352403:349392],tree_6[231923:228912],tree_6[234935:231924]);
csa_3012 csau_3012_i1346(tree_5[355415:352404],tree_5[358427:355416],tree_5[361439:358428],tree_6[237947:234936],tree_6[240959:237948]);
csa_3012 csau_3012_i1347(tree_5[364451:361440],tree_5[367463:364452],tree_5[370475:367464],tree_6[243971:240960],tree_6[246983:243972]);
csa_3012 csau_3012_i1348(tree_5[373487:370476],tree_5[376499:373488],tree_5[379511:376500],tree_6[249995:246984],tree_6[253007:249996]);
csa_3012 csau_3012_i1349(tree_5[382523:379512],tree_5[385535:382524],tree_5[388547:385536],tree_6[256019:253008],tree_6[259031:256020]);
csa_3012 csau_3012_i1350(tree_5[391559:388548],tree_5[394571:391560],tree_5[397583:394572],tree_6[262043:259032],tree_6[265055:262044]);
csa_3012 csau_3012_i1351(tree_5[400595:397584],tree_5[403607:400596],tree_5[406619:403608],tree_6[268067:265056],tree_6[271079:268068]);
csa_3012 csau_3012_i1352(tree_5[409631:406620],tree_5[412643:409632],tree_5[415655:412644],tree_6[274091:271080],tree_6[277103:274092]);
csa_3012 csau_3012_i1353(tree_5[418667:415656],tree_5[421679:418668],tree_5[424691:421680],tree_6[280115:277104],tree_6[283127:280116]);
csa_3012 csau_3012_i1354(tree_5[427703:424692],tree_5[430715:427704],tree_5[433727:430716],tree_6[286139:283128],tree_6[289151:286140]);
csa_3012 csau_3012_i1355(tree_5[436739:433728],tree_5[439751:436740],tree_5[442763:439752],tree_6[292163:289152],tree_6[295175:292164]);
csa_3012 csau_3012_i1356(tree_5[445775:442764],tree_5[448787:445776],tree_5[451799:448788],tree_6[298187:295176],tree_6[301199:298188]);
csa_3012 csau_3012_i1357(tree_5[454811:451800],tree_5[457823:454812],tree_5[460835:457824],tree_6[304211:301200],tree_6[307223:304212]);
csa_3012 csau_3012_i1358(tree_5[463847:460836],tree_5[466859:463848],tree_5[469871:466860],tree_6[310235:307224],tree_6[313247:310236]);
csa_3012 csau_3012_i1359(tree_5[472883:469872],tree_5[475895:472884],tree_5[478907:475896],tree_6[316259:313248],tree_6[319271:316260]);
csa_3012 csau_3012_i1360(tree_5[481919:478908],tree_5[484931:481920],tree_5[487943:484932],tree_6[322283:319272],tree_6[325295:322284]);
csa_3012 csau_3012_i1361(tree_5[490955:487944],tree_5[493967:490956],tree_5[496979:493968],tree_6[328307:325296],tree_6[331319:328308]);
csa_3012 csau_3012_i1362(tree_5[499991:496980],tree_5[503003:499992],tree_5[506015:503004],tree_6[334331:331320],tree_6[337343:334332]);
csa_3012 csau_3012_i1363(tree_5[509027:506016],tree_5[512039:509028],tree_5[515051:512040],tree_6[340355:337344],tree_6[343367:340356]);
csa_3012 csau_3012_i1364(tree_5[518063:515052],tree_5[521075:518064],tree_5[524087:521076],tree_6[346379:343368],tree_6[349391:346380]);
csa_3012 csau_3012_i1365(tree_5[527099:524088],tree_5[530111:527100],tree_5[533123:530112],tree_6[352403:349392],tree_6[355415:352404]);
csa_3012 csau_3012_i1366(tree_5[536135:533124],tree_5[539147:536136],tree_5[542159:539148],tree_6[358427:355416],tree_6[361439:358428]);
csa_3012 csau_3012_i1367(tree_5[545171:542160],tree_5[548183:545172],tree_5[551195:548184],tree_6[364451:361440],tree_6[367463:364452]);
csa_3012 csau_3012_i1368(tree_5[554207:551196],tree_5[557219:554208],tree_5[560231:557220],tree_6[370475:367464],tree_6[373487:370476]);
csa_3012 csau_3012_i1369(tree_5[563243:560232],tree_5[566255:563244],tree_5[569267:566256],tree_6[376499:373488],tree_6[379511:376500]);
csa_3012 csau_3012_i1370(tree_5[572279:569268],tree_5[575291:572280],tree_5[578303:575292],tree_6[382523:379512],tree_6[385535:382524]);
csa_3012 csau_3012_i1371(tree_5[581315:578304],tree_5[584327:581316],tree_5[587339:584328],tree_6[388547:385536],tree_6[391559:388548]);
csa_3012 csau_3012_i1372(tree_5[590351:587340],tree_5[593363:590352],tree_5[596375:593364],tree_6[394571:391560],tree_6[397583:394572]);
assign tree_6[400595:397584] = tree_5[599387:596376];
// layer-7
csa_3012 csau_3012_i1373(tree_6[3011:0],tree_6[6023:3012],tree_6[9035:6024],tree_7[3011:0],tree_7[6023:3012]);
csa_3012 csau_3012_i1374(tree_6[12047:9036],tree_6[15059:12048],tree_6[18071:15060],tree_7[9035:6024],tree_7[12047:9036]);
csa_3012 csau_3012_i1375(tree_6[21083:18072],tree_6[24095:21084],tree_6[27107:24096],tree_7[15059:12048],tree_7[18071:15060]);
csa_3012 csau_3012_i1376(tree_6[30119:27108],tree_6[33131:30120],tree_6[36143:33132],tree_7[21083:18072],tree_7[24095:21084]);
csa_3012 csau_3012_i1377(tree_6[39155:36144],tree_6[42167:39156],tree_6[45179:42168],tree_7[27107:24096],tree_7[30119:27108]);
csa_3012 csau_3012_i1378(tree_6[48191:45180],tree_6[51203:48192],tree_6[54215:51204],tree_7[33131:30120],tree_7[36143:33132]);
csa_3012 csau_3012_i1379(tree_6[57227:54216],tree_6[60239:57228],tree_6[63251:60240],tree_7[39155:36144],tree_7[42167:39156]);
csa_3012 csau_3012_i1380(tree_6[66263:63252],tree_6[69275:66264],tree_6[72287:69276],tree_7[45179:42168],tree_7[48191:45180]);
csa_3012 csau_3012_i1381(tree_6[75299:72288],tree_6[78311:75300],tree_6[81323:78312],tree_7[51203:48192],tree_7[54215:51204]);
csa_3012 csau_3012_i1382(tree_6[84335:81324],tree_6[87347:84336],tree_6[90359:87348],tree_7[57227:54216],tree_7[60239:57228]);
csa_3012 csau_3012_i1383(tree_6[93371:90360],tree_6[96383:93372],tree_6[99395:96384],tree_7[63251:60240],tree_7[66263:63252]);
csa_3012 csau_3012_i1384(tree_6[102407:99396],tree_6[105419:102408],tree_6[108431:105420],tree_7[69275:66264],tree_7[72287:69276]);
csa_3012 csau_3012_i1385(tree_6[111443:108432],tree_6[114455:111444],tree_6[117467:114456],tree_7[75299:72288],tree_7[78311:75300]);
csa_3012 csau_3012_i1386(tree_6[120479:117468],tree_6[123491:120480],tree_6[126503:123492],tree_7[81323:78312],tree_7[84335:81324]);
csa_3012 csau_3012_i1387(tree_6[129515:126504],tree_6[132527:129516],tree_6[135539:132528],tree_7[87347:84336],tree_7[90359:87348]);
csa_3012 csau_3012_i1388(tree_6[138551:135540],tree_6[141563:138552],tree_6[144575:141564],tree_7[93371:90360],tree_7[96383:93372]);
csa_3012 csau_3012_i1389(tree_6[147587:144576],tree_6[150599:147588],tree_6[153611:150600],tree_7[99395:96384],tree_7[102407:99396]);
csa_3012 csau_3012_i1390(tree_6[156623:153612],tree_6[159635:156624],tree_6[162647:159636],tree_7[105419:102408],tree_7[108431:105420]);
csa_3012 csau_3012_i1391(tree_6[165659:162648],tree_6[168671:165660],tree_6[171683:168672],tree_7[111443:108432],tree_7[114455:111444]);
csa_3012 csau_3012_i1392(tree_6[174695:171684],tree_6[177707:174696],tree_6[180719:177708],tree_7[117467:114456],tree_7[120479:117468]);
csa_3012 csau_3012_i1393(tree_6[183731:180720],tree_6[186743:183732],tree_6[189755:186744],tree_7[123491:120480],tree_7[126503:123492]);
csa_3012 csau_3012_i1394(tree_6[192767:189756],tree_6[195779:192768],tree_6[198791:195780],tree_7[129515:126504],tree_7[132527:129516]);
csa_3012 csau_3012_i1395(tree_6[201803:198792],tree_6[204815:201804],tree_6[207827:204816],tree_7[135539:132528],tree_7[138551:135540]);
csa_3012 csau_3012_i1396(tree_6[210839:207828],tree_6[213851:210840],tree_6[216863:213852],tree_7[141563:138552],tree_7[144575:141564]);
csa_3012 csau_3012_i1397(tree_6[219875:216864],tree_6[222887:219876],tree_6[225899:222888],tree_7[147587:144576],tree_7[150599:147588]);
csa_3012 csau_3012_i1398(tree_6[228911:225900],tree_6[231923:228912],tree_6[234935:231924],tree_7[153611:150600],tree_7[156623:153612]);
csa_3012 csau_3012_i1399(tree_6[237947:234936],tree_6[240959:237948],tree_6[243971:240960],tree_7[159635:156624],tree_7[162647:159636]);
csa_3012 csau_3012_i1400(tree_6[246983:243972],tree_6[249995:246984],tree_6[253007:249996],tree_7[165659:162648],tree_7[168671:165660]);
csa_3012 csau_3012_i1401(tree_6[256019:253008],tree_6[259031:256020],tree_6[262043:259032],tree_7[171683:168672],tree_7[174695:171684]);
csa_3012 csau_3012_i1402(tree_6[265055:262044],tree_6[268067:265056],tree_6[271079:268068],tree_7[177707:174696],tree_7[180719:177708]);
csa_3012 csau_3012_i1403(tree_6[274091:271080],tree_6[277103:274092],tree_6[280115:277104],tree_7[183731:180720],tree_7[186743:183732]);
csa_3012 csau_3012_i1404(tree_6[283127:280116],tree_6[286139:283128],tree_6[289151:286140],tree_7[189755:186744],tree_7[192767:189756]);
csa_3012 csau_3012_i1405(tree_6[292163:289152],tree_6[295175:292164],tree_6[298187:295176],tree_7[195779:192768],tree_7[198791:195780]);
csa_3012 csau_3012_i1406(tree_6[301199:298188],tree_6[304211:301200],tree_6[307223:304212],tree_7[201803:198792],tree_7[204815:201804]);
csa_3012 csau_3012_i1407(tree_6[310235:307224],tree_6[313247:310236],tree_6[316259:313248],tree_7[207827:204816],tree_7[210839:207828]);
csa_3012 csau_3012_i1408(tree_6[319271:316260],tree_6[322283:319272],tree_6[325295:322284],tree_7[213851:210840],tree_7[216863:213852]);
csa_3012 csau_3012_i1409(tree_6[328307:325296],tree_6[331319:328308],tree_6[334331:331320],tree_7[219875:216864],tree_7[222887:219876]);
csa_3012 csau_3012_i1410(tree_6[337343:334332],tree_6[340355:337344],tree_6[343367:340356],tree_7[225899:222888],tree_7[228911:225900]);
csa_3012 csau_3012_i1411(tree_6[346379:343368],tree_6[349391:346380],tree_6[352403:349392],tree_7[231923:228912],tree_7[234935:231924]);
csa_3012 csau_3012_i1412(tree_6[355415:352404],tree_6[358427:355416],tree_6[361439:358428],tree_7[237947:234936],tree_7[240959:237948]);
csa_3012 csau_3012_i1413(tree_6[364451:361440],tree_6[367463:364452],tree_6[370475:367464],tree_7[243971:240960],tree_7[246983:243972]);
csa_3012 csau_3012_i1414(tree_6[373487:370476],tree_6[376499:373488],tree_6[379511:376500],tree_7[249995:246984],tree_7[253007:249996]);
csa_3012 csau_3012_i1415(tree_6[382523:379512],tree_6[385535:382524],tree_6[388547:385536],tree_7[256019:253008],tree_7[259031:256020]);
csa_3012 csau_3012_i1416(tree_6[391559:388548],tree_6[394571:391560],tree_6[397583:394572],tree_7[262043:259032],tree_7[265055:262044]);
assign tree_7[268067:265056] = tree_6[400595:397584];
// layer-8
csa_3012 csau_3012_i1417(tree_7[3011:0],tree_7[6023:3012],tree_7[9035:6024],tree_8[3011:0],tree_8[6023:3012]);
csa_3012 csau_3012_i1418(tree_7[12047:9036],tree_7[15059:12048],tree_7[18071:15060],tree_8[9035:6024],tree_8[12047:9036]);
csa_3012 csau_3012_i1419(tree_7[21083:18072],tree_7[24095:21084],tree_7[27107:24096],tree_8[15059:12048],tree_8[18071:15060]);
csa_3012 csau_3012_i1420(tree_7[30119:27108],tree_7[33131:30120],tree_7[36143:33132],tree_8[21083:18072],tree_8[24095:21084]);
csa_3012 csau_3012_i1421(tree_7[39155:36144],tree_7[42167:39156],tree_7[45179:42168],tree_8[27107:24096],tree_8[30119:27108]);
csa_3012 csau_3012_i1422(tree_7[48191:45180],tree_7[51203:48192],tree_7[54215:51204],tree_8[33131:30120],tree_8[36143:33132]);
csa_3012 csau_3012_i1423(tree_7[57227:54216],tree_7[60239:57228],tree_7[63251:60240],tree_8[39155:36144],tree_8[42167:39156]);
csa_3012 csau_3012_i1424(tree_7[66263:63252],tree_7[69275:66264],tree_7[72287:69276],tree_8[45179:42168],tree_8[48191:45180]);
csa_3012 csau_3012_i1425(tree_7[75299:72288],tree_7[78311:75300],tree_7[81323:78312],tree_8[51203:48192],tree_8[54215:51204]);
csa_3012 csau_3012_i1426(tree_7[84335:81324],tree_7[87347:84336],tree_7[90359:87348],tree_8[57227:54216],tree_8[60239:57228]);
csa_3012 csau_3012_i1427(tree_7[93371:90360],tree_7[96383:93372],tree_7[99395:96384],tree_8[63251:60240],tree_8[66263:63252]);
csa_3012 csau_3012_i1428(tree_7[102407:99396],tree_7[105419:102408],tree_7[108431:105420],tree_8[69275:66264],tree_8[72287:69276]);
csa_3012 csau_3012_i1429(tree_7[111443:108432],tree_7[114455:111444],tree_7[117467:114456],tree_8[75299:72288],tree_8[78311:75300]);
csa_3012 csau_3012_i1430(tree_7[120479:117468],tree_7[123491:120480],tree_7[126503:123492],tree_8[81323:78312],tree_8[84335:81324]);
csa_3012 csau_3012_i1431(tree_7[129515:126504],tree_7[132527:129516],tree_7[135539:132528],tree_8[87347:84336],tree_8[90359:87348]);
csa_3012 csau_3012_i1432(tree_7[138551:135540],tree_7[141563:138552],tree_7[144575:141564],tree_8[93371:90360],tree_8[96383:93372]);
csa_3012 csau_3012_i1433(tree_7[147587:144576],tree_7[150599:147588],tree_7[153611:150600],tree_8[99395:96384],tree_8[102407:99396]);
csa_3012 csau_3012_i1434(tree_7[156623:153612],tree_7[159635:156624],tree_7[162647:159636],tree_8[105419:102408],tree_8[108431:105420]);
csa_3012 csau_3012_i1435(tree_7[165659:162648],tree_7[168671:165660],tree_7[171683:168672],tree_8[111443:108432],tree_8[114455:111444]);
csa_3012 csau_3012_i1436(tree_7[174695:171684],tree_7[177707:174696],tree_7[180719:177708],tree_8[117467:114456],tree_8[120479:117468]);
csa_3012 csau_3012_i1437(tree_7[183731:180720],tree_7[186743:183732],tree_7[189755:186744],tree_8[123491:120480],tree_8[126503:123492]);
csa_3012 csau_3012_i1438(tree_7[192767:189756],tree_7[195779:192768],tree_7[198791:195780],tree_8[129515:126504],tree_8[132527:129516]);
csa_3012 csau_3012_i1439(tree_7[201803:198792],tree_7[204815:201804],tree_7[207827:204816],tree_8[135539:132528],tree_8[138551:135540]);
csa_3012 csau_3012_i1440(tree_7[210839:207828],tree_7[213851:210840],tree_7[216863:213852],tree_8[141563:138552],tree_8[144575:141564]);
csa_3012 csau_3012_i1441(tree_7[219875:216864],tree_7[222887:219876],tree_7[225899:222888],tree_8[147587:144576],tree_8[150599:147588]);
csa_3012 csau_3012_i1442(tree_7[228911:225900],tree_7[231923:228912],tree_7[234935:231924],tree_8[153611:150600],tree_8[156623:153612]);
csa_3012 csau_3012_i1443(tree_7[237947:234936],tree_7[240959:237948],tree_7[243971:240960],tree_8[159635:156624],tree_8[162647:159636]);
csa_3012 csau_3012_i1444(tree_7[246983:243972],tree_7[249995:246984],tree_7[253007:249996],tree_8[165659:162648],tree_8[168671:165660]);
csa_3012 csau_3012_i1445(tree_7[256019:253008],tree_7[259031:256020],tree_7[262043:259032],tree_8[171683:168672],tree_8[174695:171684]);
assign tree_8[177707:174696] = tree_7[265055:262044];
assign tree_8[180719:177708] = tree_7[268067:265056];
// layer-9
csa_3012 csau_3012_i1446(tree_8[3011:0],tree_8[6023:3012],tree_8[9035:6024],tree_9[3011:0],tree_9[6023:3012]);
csa_3012 csau_3012_i1447(tree_8[12047:9036],tree_8[15059:12048],tree_8[18071:15060],tree_9[9035:6024],tree_9[12047:9036]);
csa_3012 csau_3012_i1448(tree_8[21083:18072],tree_8[24095:21084],tree_8[27107:24096],tree_9[15059:12048],tree_9[18071:15060]);
csa_3012 csau_3012_i1449(tree_8[30119:27108],tree_8[33131:30120],tree_8[36143:33132],tree_9[21083:18072],tree_9[24095:21084]);
csa_3012 csau_3012_i1450(tree_8[39155:36144],tree_8[42167:39156],tree_8[45179:42168],tree_9[27107:24096],tree_9[30119:27108]);
csa_3012 csau_3012_i1451(tree_8[48191:45180],tree_8[51203:48192],tree_8[54215:51204],tree_9[33131:30120],tree_9[36143:33132]);
csa_3012 csau_3012_i1452(tree_8[57227:54216],tree_8[60239:57228],tree_8[63251:60240],tree_9[39155:36144],tree_9[42167:39156]);
csa_3012 csau_3012_i1453(tree_8[66263:63252],tree_8[69275:66264],tree_8[72287:69276],tree_9[45179:42168],tree_9[48191:45180]);
csa_3012 csau_3012_i1454(tree_8[75299:72288],tree_8[78311:75300],tree_8[81323:78312],tree_9[51203:48192],tree_9[54215:51204]);
csa_3012 csau_3012_i1455(tree_8[84335:81324],tree_8[87347:84336],tree_8[90359:87348],tree_9[57227:54216],tree_9[60239:57228]);
csa_3012 csau_3012_i1456(tree_8[93371:90360],tree_8[96383:93372],tree_8[99395:96384],tree_9[63251:60240],tree_9[66263:63252]);
csa_3012 csau_3012_i1457(tree_8[102407:99396],tree_8[105419:102408],tree_8[108431:105420],tree_9[69275:66264],tree_9[72287:69276]);
csa_3012 csau_3012_i1458(tree_8[111443:108432],tree_8[114455:111444],tree_8[117467:114456],tree_9[75299:72288],tree_9[78311:75300]);
csa_3012 csau_3012_i1459(tree_8[120479:117468],tree_8[123491:120480],tree_8[126503:123492],tree_9[81323:78312],tree_9[84335:81324]);
csa_3012 csau_3012_i1460(tree_8[129515:126504],tree_8[132527:129516],tree_8[135539:132528],tree_9[87347:84336],tree_9[90359:87348]);
csa_3012 csau_3012_i1461(tree_8[138551:135540],tree_8[141563:138552],tree_8[144575:141564],tree_9[93371:90360],tree_9[96383:93372]);
csa_3012 csau_3012_i1462(tree_8[147587:144576],tree_8[150599:147588],tree_8[153611:150600],tree_9[99395:96384],tree_9[102407:99396]);
csa_3012 csau_3012_i1463(tree_8[156623:153612],tree_8[159635:156624],tree_8[162647:159636],tree_9[105419:102408],tree_9[108431:105420]);
csa_3012 csau_3012_i1464(tree_8[165659:162648],tree_8[168671:165660],tree_8[171683:168672],tree_9[111443:108432],tree_9[114455:111444]);
csa_3012 csau_3012_i1465(tree_8[174695:171684],tree_8[177707:174696],tree_8[180719:177708],tree_9[117467:114456],tree_9[120479:117468]);
// layer-10
csa_3012 csau_3012_i1466(tree_9[3011:0],tree_9[6023:3012],tree_9[9035:6024],tree_10[3011:0],tree_10[6023:3012]);
csa_3012 csau_3012_i1467(tree_9[12047:9036],tree_9[15059:12048],tree_9[18071:15060],tree_10[9035:6024],tree_10[12047:9036]);
csa_3012 csau_3012_i1468(tree_9[21083:18072],tree_9[24095:21084],tree_9[27107:24096],tree_10[15059:12048],tree_10[18071:15060]);
csa_3012 csau_3012_i1469(tree_9[30119:27108],tree_9[33131:30120],tree_9[36143:33132],tree_10[21083:18072],tree_10[24095:21084]);
csa_3012 csau_3012_i1470(tree_9[39155:36144],tree_9[42167:39156],tree_9[45179:42168],tree_10[27107:24096],tree_10[30119:27108]);
csa_3012 csau_3012_i1471(tree_9[48191:45180],tree_9[51203:48192],tree_9[54215:51204],tree_10[33131:30120],tree_10[36143:33132]);
csa_3012 csau_3012_i1472(tree_9[57227:54216],tree_9[60239:57228],tree_9[63251:60240],tree_10[39155:36144],tree_10[42167:39156]);
csa_3012 csau_3012_i1473(tree_9[66263:63252],tree_9[69275:66264],tree_9[72287:69276],tree_10[45179:42168],tree_10[48191:45180]);
csa_3012 csau_3012_i1474(tree_9[75299:72288],tree_9[78311:75300],tree_9[81323:78312],tree_10[51203:48192],tree_10[54215:51204]);
csa_3012 csau_3012_i1475(tree_9[84335:81324],tree_9[87347:84336],tree_9[90359:87348],tree_10[57227:54216],tree_10[60239:57228]);
csa_3012 csau_3012_i1476(tree_9[93371:90360],tree_9[96383:93372],tree_9[99395:96384],tree_10[63251:60240],tree_10[66263:63252]);
csa_3012 csau_3012_i1477(tree_9[102407:99396],tree_9[105419:102408],tree_9[108431:105420],tree_10[69275:66264],tree_10[72287:69276]);
csa_3012 csau_3012_i1478(tree_9[111443:108432],tree_9[114455:111444],tree_9[117467:114456],tree_10[75299:72288],tree_10[78311:75300]);
assign tree_10[81323:78312] = tree_9[120479:117468];
// layer-11
csa_3012 csau_3012_i1479(tree_10[3011:0],tree_10[6023:3012],tree_10[9035:6024],tree_11[3011:0],tree_11[6023:3012]);
csa_3012 csau_3012_i1480(tree_10[12047:9036],tree_10[15059:12048],tree_10[18071:15060],tree_11[9035:6024],tree_11[12047:9036]);
csa_3012 csau_3012_i1481(tree_10[21083:18072],tree_10[24095:21084],tree_10[27107:24096],tree_11[15059:12048],tree_11[18071:15060]);
csa_3012 csau_3012_i1482(tree_10[30119:27108],tree_10[33131:30120],tree_10[36143:33132],tree_11[21083:18072],tree_11[24095:21084]);
csa_3012 csau_3012_i1483(tree_10[39155:36144],tree_10[42167:39156],tree_10[45179:42168],tree_11[27107:24096],tree_11[30119:27108]);
csa_3012 csau_3012_i1484(tree_10[48191:45180],tree_10[51203:48192],tree_10[54215:51204],tree_11[33131:30120],tree_11[36143:33132]);
csa_3012 csau_3012_i1485(tree_10[57227:54216],tree_10[60239:57228],tree_10[63251:60240],tree_11[39155:36144],tree_11[42167:39156]);
csa_3012 csau_3012_i1486(tree_10[66263:63252],tree_10[69275:66264],tree_10[72287:69276],tree_11[45179:42168],tree_11[48191:45180]);
csa_3012 csau_3012_i1487(tree_10[75299:72288],tree_10[78311:75300],tree_10[81323:78312],tree_11[51203:48192],tree_11[54215:51204]);
// layer-12
csa_3012 csau_3012_i1488(tree_11[3011:0],tree_11[6023:3012],tree_11[9035:6024],tree_12[3011:0],tree_12[6023:3012]);
csa_3012 csau_3012_i1489(tree_11[12047:9036],tree_11[15059:12048],tree_11[18071:15060],tree_12[9035:6024],tree_12[12047:9036]);
csa_3012 csau_3012_i1490(tree_11[21083:18072],tree_11[24095:21084],tree_11[27107:24096],tree_12[15059:12048],tree_12[18071:15060]);
csa_3012 csau_3012_i1491(tree_11[30119:27108],tree_11[33131:30120],tree_11[36143:33132],tree_12[21083:18072],tree_12[24095:21084]);
csa_3012 csau_3012_i1492(tree_11[39155:36144],tree_11[42167:39156],tree_11[45179:42168],tree_12[27107:24096],tree_12[30119:27108]);
csa_3012 csau_3012_i1493(tree_11[48191:45180],tree_11[51203:48192],tree_11[54215:51204],tree_12[33131:30120],tree_12[36143:33132]);
// layer-13
csa_3012 csau_3012_i1494(tree_12[3011:0],tree_12[6023:3012],tree_12[9035:6024],tree_13[3011:0],tree_13[6023:3012]);
csa_3012 csau_3012_i1495(tree_12[12047:9036],tree_12[15059:12048],tree_12[18071:15060],tree_13[9035:6024],tree_13[12047:9036]);
csa_3012 csau_3012_i1496(tree_12[21083:18072],tree_12[24095:21084],tree_12[27107:24096],tree_13[15059:12048],tree_13[18071:15060]);
csa_3012 csau_3012_i1497(tree_12[30119:27108],tree_12[33131:30120],tree_12[36143:33132],tree_13[21083:18072],tree_13[24095:21084]);
// layer-14
csa_3012 csau_3012_i1498(tree_13[3011:0],tree_13[6023:3012],tree_13[9035:6024],tree_14[3011:0],tree_14[6023:3012]);
csa_3012 csau_3012_i1499(tree_13[12047:9036],tree_13[15059:12048],tree_13[18071:15060],tree_14[9035:6024],tree_14[12047:9036]);
assign tree_14[15059:12048] = tree_13[21083:18072];
assign tree_14[18071:15060] = tree_13[24095:21084];
// layer-15
csa_3012 csau_3012_i1500(tree_14[3011:0],tree_14[6023:3012],tree_14[9035:6024],tree_15[3011:0],tree_15[6023:3012]);
csa_3012 csau_3012_i1501(tree_14[12047:9036],tree_14[15059:12048],tree_14[18071:15060],tree_15[9035:6024],tree_15[12047:9036]);
// layer-16
csa_3012 csau_3012_i1502(tree_15[3011:0],tree_15[6023:3012],tree_15[9035:6024],tree_16[3011:0],tree_16[6023:3012]);
assign tree_16[9035:6024] = tree_15[12047:9036];
// layer-17
csa_3012 csau_3012_i1503(tree_16[3011:0],tree_16[6023:3012],tree_16[9035:6024],tree_17[3011:0],tree_17[6023:3012]);

// final assignment
assign B_0 = tree_17[3011:0];
assign B_1 = tree_17[6023:3012];

endmodule
