

module csa_tree_92x92_truncated(
    input [8463:0] A, // lines are appended together
    output[91:0] B_0,
    output[91:0] B_1
);

wire [5703:0] tree_1;
wire [3863:0] tree_2;
wire [2575:0] tree_3;
wire [1747:0] tree_4;
wire [1195:0] tree_5;
wire [827:0] tree_6;
wire [551:0] tree_7;
wire [367:0] tree_8;
wire [275:0] tree_9;
wire [183:0] tree_10;
// layer-1
csa_92 csau_92_i0(A[91:0],A[183:92],A[275:184],tree_1[91:0],tree_1[183:92]);
csa_92 csau_92_i1(A[367:276],A[459:368],A[551:460],tree_1[275:184],tree_1[367:276]);
csa_92 csau_92_i2(A[643:552],A[735:644],A[827:736],tree_1[459:368],tree_1[551:460]);
csa_92 csau_92_i3(A[919:828],A[1011:920],A[1103:1012],tree_1[643:552],tree_1[735:644]);
csa_92 csau_92_i4(A[1195:1104],A[1287:1196],A[1379:1288],tree_1[827:736],tree_1[919:828]);
csa_92 csau_92_i5(A[1471:1380],A[1563:1472],A[1655:1564],tree_1[1011:920],tree_1[1103:1012]);
csa_92 csau_92_i6(A[1747:1656],A[1839:1748],A[1931:1840],tree_1[1195:1104],tree_1[1287:1196]);
csa_92 csau_92_i7(A[2023:1932],A[2115:2024],A[2207:2116],tree_1[1379:1288],tree_1[1471:1380]);
csa_92 csau_92_i8(A[2299:2208],A[2391:2300],A[2483:2392],tree_1[1563:1472],tree_1[1655:1564]);
csa_92 csau_92_i9(A[2575:2484],A[2667:2576],A[2759:2668],tree_1[1747:1656],tree_1[1839:1748]);
csa_92 csau_92_i10(A[2851:2760],A[2943:2852],A[3035:2944],tree_1[1931:1840],tree_1[2023:1932]);
csa_92 csau_92_i11(A[3127:3036],A[3219:3128],A[3311:3220],tree_1[2115:2024],tree_1[2207:2116]);
csa_92 csau_92_i12(A[3403:3312],A[3495:3404],A[3587:3496],tree_1[2299:2208],tree_1[2391:2300]);
csa_92 csau_92_i13(A[3679:3588],A[3771:3680],A[3863:3772],tree_1[2483:2392],tree_1[2575:2484]);
csa_92 csau_92_i14(A[3955:3864],A[4047:3956],A[4139:4048],tree_1[2667:2576],tree_1[2759:2668]);
csa_92 csau_92_i15(A[4231:4140],A[4323:4232],A[4415:4324],tree_1[2851:2760],tree_1[2943:2852]);
csa_92 csau_92_i16(A[4507:4416],A[4599:4508],A[4691:4600],tree_1[3035:2944],tree_1[3127:3036]);
csa_92 csau_92_i17(A[4783:4692],A[4875:4784],A[4967:4876],tree_1[3219:3128],tree_1[3311:3220]);
csa_92 csau_92_i18(A[5059:4968],A[5151:5060],A[5243:5152],tree_1[3403:3312],tree_1[3495:3404]);
csa_92 csau_92_i19(A[5335:5244],A[5427:5336],A[5519:5428],tree_1[3587:3496],tree_1[3679:3588]);
csa_92 csau_92_i20(A[5611:5520],A[5703:5612],A[5795:5704],tree_1[3771:3680],tree_1[3863:3772]);
csa_92 csau_92_i21(A[5887:5796],A[5979:5888],A[6071:5980],tree_1[3955:3864],tree_1[4047:3956]);
csa_92 csau_92_i22(A[6163:6072],A[6255:6164],A[6347:6256],tree_1[4139:4048],tree_1[4231:4140]);
csa_92 csau_92_i23(A[6439:6348],A[6531:6440],A[6623:6532],tree_1[4323:4232],tree_1[4415:4324]);
csa_92 csau_92_i24(A[6715:6624],A[6807:6716],A[6899:6808],tree_1[4507:4416],tree_1[4599:4508]);
csa_92 csau_92_i25(A[6991:6900],A[7083:6992],A[7175:7084],tree_1[4691:4600],tree_1[4783:4692]);
csa_92 csau_92_i26(A[7267:7176],A[7359:7268],A[7451:7360],tree_1[4875:4784],tree_1[4967:4876]);
csa_92 csau_92_i27(A[7543:7452],A[7635:7544],A[7727:7636],tree_1[5059:4968],tree_1[5151:5060]);
csa_92 csau_92_i28(A[7819:7728],A[7911:7820],A[8003:7912],tree_1[5243:5152],tree_1[5335:5244]);
csa_92 csau_92_i29(A[8095:8004],A[8187:8096],A[8279:8188],tree_1[5427:5336],tree_1[5519:5428]);
assign tree_1[5611:5520] = A[8371:8280];
assign tree_1[5703:5612] = A[8463:8372];
// layer-2
csa_92 csau_92_i30(tree_1[91:0],tree_1[183:92],tree_1[275:184],tree_2[91:0],tree_2[183:92]);
csa_92 csau_92_i31(tree_1[367:276],tree_1[459:368],tree_1[551:460],tree_2[275:184],tree_2[367:276]);
csa_92 csau_92_i32(tree_1[643:552],tree_1[735:644],tree_1[827:736],tree_2[459:368],tree_2[551:460]);
csa_92 csau_92_i33(tree_1[919:828],tree_1[1011:920],tree_1[1103:1012],tree_2[643:552],tree_2[735:644]);
csa_92 csau_92_i34(tree_1[1195:1104],tree_1[1287:1196],tree_1[1379:1288],tree_2[827:736],tree_2[919:828]);
csa_92 csau_92_i35(tree_1[1471:1380],tree_1[1563:1472],tree_1[1655:1564],tree_2[1011:920],tree_2[1103:1012]);
csa_92 csau_92_i36(tree_1[1747:1656],tree_1[1839:1748],tree_1[1931:1840],tree_2[1195:1104],tree_2[1287:1196]);
csa_92 csau_92_i37(tree_1[2023:1932],tree_1[2115:2024],tree_1[2207:2116],tree_2[1379:1288],tree_2[1471:1380]);
csa_92 csau_92_i38(tree_1[2299:2208],tree_1[2391:2300],tree_1[2483:2392],tree_2[1563:1472],tree_2[1655:1564]);
csa_92 csau_92_i39(tree_1[2575:2484],tree_1[2667:2576],tree_1[2759:2668],tree_2[1747:1656],tree_2[1839:1748]);
csa_92 csau_92_i40(tree_1[2851:2760],tree_1[2943:2852],tree_1[3035:2944],tree_2[1931:1840],tree_2[2023:1932]);
csa_92 csau_92_i41(tree_1[3127:3036],tree_1[3219:3128],tree_1[3311:3220],tree_2[2115:2024],tree_2[2207:2116]);
csa_92 csau_92_i42(tree_1[3403:3312],tree_1[3495:3404],tree_1[3587:3496],tree_2[2299:2208],tree_2[2391:2300]);
csa_92 csau_92_i43(tree_1[3679:3588],tree_1[3771:3680],tree_1[3863:3772],tree_2[2483:2392],tree_2[2575:2484]);
csa_92 csau_92_i44(tree_1[3955:3864],tree_1[4047:3956],tree_1[4139:4048],tree_2[2667:2576],tree_2[2759:2668]);
csa_92 csau_92_i45(tree_1[4231:4140],tree_1[4323:4232],tree_1[4415:4324],tree_2[2851:2760],tree_2[2943:2852]);
csa_92 csau_92_i46(tree_1[4507:4416],tree_1[4599:4508],tree_1[4691:4600],tree_2[3035:2944],tree_2[3127:3036]);
csa_92 csau_92_i47(tree_1[4783:4692],tree_1[4875:4784],tree_1[4967:4876],tree_2[3219:3128],tree_2[3311:3220]);
csa_92 csau_92_i48(tree_1[5059:4968],tree_1[5151:5060],tree_1[5243:5152],tree_2[3403:3312],tree_2[3495:3404]);
csa_92 csau_92_i49(tree_1[5335:5244],tree_1[5427:5336],tree_1[5519:5428],tree_2[3587:3496],tree_2[3679:3588]);
assign tree_2[3771:3680] = tree_1[5611:5520];
assign tree_2[3863:3772] = tree_1[5703:5612];
// layer-3
csa_92 csau_92_i50(tree_2[91:0],tree_2[183:92],tree_2[275:184],tree_3[91:0],tree_3[183:92]);
csa_92 csau_92_i51(tree_2[367:276],tree_2[459:368],tree_2[551:460],tree_3[275:184],tree_3[367:276]);
csa_92 csau_92_i52(tree_2[643:552],tree_2[735:644],tree_2[827:736],tree_3[459:368],tree_3[551:460]);
csa_92 csau_92_i53(tree_2[919:828],tree_2[1011:920],tree_2[1103:1012],tree_3[643:552],tree_3[735:644]);
csa_92 csau_92_i54(tree_2[1195:1104],tree_2[1287:1196],tree_2[1379:1288],tree_3[827:736],tree_3[919:828]);
csa_92 csau_92_i55(tree_2[1471:1380],tree_2[1563:1472],tree_2[1655:1564],tree_3[1011:920],tree_3[1103:1012]);
csa_92 csau_92_i56(tree_2[1747:1656],tree_2[1839:1748],tree_2[1931:1840],tree_3[1195:1104],tree_3[1287:1196]);
csa_92 csau_92_i57(tree_2[2023:1932],tree_2[2115:2024],tree_2[2207:2116],tree_3[1379:1288],tree_3[1471:1380]);
csa_92 csau_92_i58(tree_2[2299:2208],tree_2[2391:2300],tree_2[2483:2392],tree_3[1563:1472],tree_3[1655:1564]);
csa_92 csau_92_i59(tree_2[2575:2484],tree_2[2667:2576],tree_2[2759:2668],tree_3[1747:1656],tree_3[1839:1748]);
csa_92 csau_92_i60(tree_2[2851:2760],tree_2[2943:2852],tree_2[3035:2944],tree_3[1931:1840],tree_3[2023:1932]);
csa_92 csau_92_i61(tree_2[3127:3036],tree_2[3219:3128],tree_2[3311:3220],tree_3[2115:2024],tree_3[2207:2116]);
csa_92 csau_92_i62(tree_2[3403:3312],tree_2[3495:3404],tree_2[3587:3496],tree_3[2299:2208],tree_3[2391:2300]);
csa_92 csau_92_i63(tree_2[3679:3588],tree_2[3771:3680],tree_2[3863:3772],tree_3[2483:2392],tree_3[2575:2484]);
// layer-4
csa_92 csau_92_i64(tree_3[91:0],tree_3[183:92],tree_3[275:184],tree_4[91:0],tree_4[183:92]);
csa_92 csau_92_i65(tree_3[367:276],tree_3[459:368],tree_3[551:460],tree_4[275:184],tree_4[367:276]);
csa_92 csau_92_i66(tree_3[643:552],tree_3[735:644],tree_3[827:736],tree_4[459:368],tree_4[551:460]);
csa_92 csau_92_i67(tree_3[919:828],tree_3[1011:920],tree_3[1103:1012],tree_4[643:552],tree_4[735:644]);
csa_92 csau_92_i68(tree_3[1195:1104],tree_3[1287:1196],tree_3[1379:1288],tree_4[827:736],tree_4[919:828]);
csa_92 csau_92_i69(tree_3[1471:1380],tree_3[1563:1472],tree_3[1655:1564],tree_4[1011:920],tree_4[1103:1012]);
csa_92 csau_92_i70(tree_3[1747:1656],tree_3[1839:1748],tree_3[1931:1840],tree_4[1195:1104],tree_4[1287:1196]);
csa_92 csau_92_i71(tree_3[2023:1932],tree_3[2115:2024],tree_3[2207:2116],tree_4[1379:1288],tree_4[1471:1380]);
csa_92 csau_92_i72(tree_3[2299:2208],tree_3[2391:2300],tree_3[2483:2392],tree_4[1563:1472],tree_4[1655:1564]);
assign tree_4[1747:1656] = tree_3[2575:2484];
// layer-5
csa_92 csau_92_i73(tree_4[91:0],tree_4[183:92],tree_4[275:184],tree_5[91:0],tree_5[183:92]);
csa_92 csau_92_i74(tree_4[367:276],tree_4[459:368],tree_4[551:460],tree_5[275:184],tree_5[367:276]);
csa_92 csau_92_i75(tree_4[643:552],tree_4[735:644],tree_4[827:736],tree_5[459:368],tree_5[551:460]);
csa_92 csau_92_i76(tree_4[919:828],tree_4[1011:920],tree_4[1103:1012],tree_5[643:552],tree_5[735:644]);
csa_92 csau_92_i77(tree_4[1195:1104],tree_4[1287:1196],tree_4[1379:1288],tree_5[827:736],tree_5[919:828]);
csa_92 csau_92_i78(tree_4[1471:1380],tree_4[1563:1472],tree_4[1655:1564],tree_5[1011:920],tree_5[1103:1012]);
assign tree_5[1195:1104] = tree_4[1747:1656];
// layer-6
csa_92 csau_92_i79(tree_5[91:0],tree_5[183:92],tree_5[275:184],tree_6[91:0],tree_6[183:92]);
csa_92 csau_92_i80(tree_5[367:276],tree_5[459:368],tree_5[551:460],tree_6[275:184],tree_6[367:276]);
csa_92 csau_92_i81(tree_5[643:552],tree_5[735:644],tree_5[827:736],tree_6[459:368],tree_6[551:460]);
csa_92 csau_92_i82(tree_5[919:828],tree_5[1011:920],tree_5[1103:1012],tree_6[643:552],tree_6[735:644]);
assign tree_6[827:736] = tree_5[1195:1104];
// layer-7
csa_92 csau_92_i83(tree_6[91:0],tree_6[183:92],tree_6[275:184],tree_7[91:0],tree_7[183:92]);
csa_92 csau_92_i84(tree_6[367:276],tree_6[459:368],tree_6[551:460],tree_7[275:184],tree_7[367:276]);
csa_92 csau_92_i85(tree_6[643:552],tree_6[735:644],tree_6[827:736],tree_7[459:368],tree_7[551:460]);
// layer-8
csa_92 csau_92_i86(tree_7[91:0],tree_7[183:92],tree_7[275:184],tree_8[91:0],tree_8[183:92]);
csa_92 csau_92_i87(tree_7[367:276],tree_7[459:368],tree_7[551:460],tree_8[275:184],tree_8[367:276]);
// layer-9
csa_92 csau_92_i88(tree_8[91:0],tree_8[183:92],tree_8[275:184],tree_9[91:0],tree_9[183:92]);
assign tree_9[275:184] = tree_8[367:276];
// layer-10
csa_92 csau_92_i89(tree_9[91:0],tree_9[183:92],tree_9[275:184],tree_10[91:0],tree_10[183:92]);

// final assignment
assign B_0 = tree_10[91:0];
assign B_1 = tree_10[183:92];

endmodule
