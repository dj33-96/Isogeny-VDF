
module AND_matrix_1506x1506(
    input [1505:0] a,
    input [1505:0] b,
    output [4536071:0] c // lines are appended together
);
    
wire [1505:0] c_w_0;
wire [1505:0] c_w_1;
wire [1505:0] c_w_2;
wire [1505:0] c_w_3;
wire [1505:0] c_w_4;
wire [1505:0] c_w_5;
wire [1505:0] c_w_6;
wire [1505:0] c_w_7;
wire [1505:0] c_w_8;
wire [1505:0] c_w_9;
wire [1505:0] c_w_10;
wire [1505:0] c_w_11;
wire [1505:0] c_w_12;
wire [1505:0] c_w_13;
wire [1505:0] c_w_14;
wire [1505:0] c_w_15;
wire [1505:0] c_w_16;
wire [1505:0] c_w_17;
wire [1505:0] c_w_18;
wire [1505:0] c_w_19;
wire [1505:0] c_w_20;
wire [1505:0] c_w_21;
wire [1505:0] c_w_22;
wire [1505:0] c_w_23;
wire [1505:0] c_w_24;
wire [1505:0] c_w_25;
wire [1505:0] c_w_26;
wire [1505:0] c_w_27;
wire [1505:0] c_w_28;
wire [1505:0] c_w_29;
wire [1505:0] c_w_30;
wire [1505:0] c_w_31;
wire [1505:0] c_w_32;
wire [1505:0] c_w_33;
wire [1505:0] c_w_34;
wire [1505:0] c_w_35;
wire [1505:0] c_w_36;
wire [1505:0] c_w_37;
wire [1505:0] c_w_38;
wire [1505:0] c_w_39;
wire [1505:0] c_w_40;
wire [1505:0] c_w_41;
wire [1505:0] c_w_42;
wire [1505:0] c_w_43;
wire [1505:0] c_w_44;
wire [1505:0] c_w_45;
wire [1505:0] c_w_46;
wire [1505:0] c_w_47;
wire [1505:0] c_w_48;
wire [1505:0] c_w_49;
wire [1505:0] c_w_50;
wire [1505:0] c_w_51;
wire [1505:0] c_w_52;
wire [1505:0] c_w_53;
wire [1505:0] c_w_54;
wire [1505:0] c_w_55;
wire [1505:0] c_w_56;
wire [1505:0] c_w_57;
wire [1505:0] c_w_58;
wire [1505:0] c_w_59;
wire [1505:0] c_w_60;
wire [1505:0] c_w_61;
wire [1505:0] c_w_62;
wire [1505:0] c_w_63;
wire [1505:0] c_w_64;
wire [1505:0] c_w_65;
wire [1505:0] c_w_66;
wire [1505:0] c_w_67;
wire [1505:0] c_w_68;
wire [1505:0] c_w_69;
wire [1505:0] c_w_70;
wire [1505:0] c_w_71;
wire [1505:0] c_w_72;
wire [1505:0] c_w_73;
wire [1505:0] c_w_74;
wire [1505:0] c_w_75;
wire [1505:0] c_w_76;
wire [1505:0] c_w_77;
wire [1505:0] c_w_78;
wire [1505:0] c_w_79;
wire [1505:0] c_w_80;
wire [1505:0] c_w_81;
wire [1505:0] c_w_82;
wire [1505:0] c_w_83;
wire [1505:0] c_w_84;
wire [1505:0] c_w_85;
wire [1505:0] c_w_86;
wire [1505:0] c_w_87;
wire [1505:0] c_w_88;
wire [1505:0] c_w_89;
wire [1505:0] c_w_90;
wire [1505:0] c_w_91;
wire [1505:0] c_w_92;
wire [1505:0] c_w_93;
wire [1505:0] c_w_94;
wire [1505:0] c_w_95;
wire [1505:0] c_w_96;
wire [1505:0] c_w_97;
wire [1505:0] c_w_98;
wire [1505:0] c_w_99;
wire [1505:0] c_w_100;
wire [1505:0] c_w_101;
wire [1505:0] c_w_102;
wire [1505:0] c_w_103;
wire [1505:0] c_w_104;
wire [1505:0] c_w_105;
wire [1505:0] c_w_106;
wire [1505:0] c_w_107;
wire [1505:0] c_w_108;
wire [1505:0] c_w_109;
wire [1505:0] c_w_110;
wire [1505:0] c_w_111;
wire [1505:0] c_w_112;
wire [1505:0] c_w_113;
wire [1505:0] c_w_114;
wire [1505:0] c_w_115;
wire [1505:0] c_w_116;
wire [1505:0] c_w_117;
wire [1505:0] c_w_118;
wire [1505:0] c_w_119;
wire [1505:0] c_w_120;
wire [1505:0] c_w_121;
wire [1505:0] c_w_122;
wire [1505:0] c_w_123;
wire [1505:0] c_w_124;
wire [1505:0] c_w_125;
wire [1505:0] c_w_126;
wire [1505:0] c_w_127;
wire [1505:0] c_w_128;
wire [1505:0] c_w_129;
wire [1505:0] c_w_130;
wire [1505:0] c_w_131;
wire [1505:0] c_w_132;
wire [1505:0] c_w_133;
wire [1505:0] c_w_134;
wire [1505:0] c_w_135;
wire [1505:0] c_w_136;
wire [1505:0] c_w_137;
wire [1505:0] c_w_138;
wire [1505:0] c_w_139;
wire [1505:0] c_w_140;
wire [1505:0] c_w_141;
wire [1505:0] c_w_142;
wire [1505:0] c_w_143;
wire [1505:0] c_w_144;
wire [1505:0] c_w_145;
wire [1505:0] c_w_146;
wire [1505:0] c_w_147;
wire [1505:0] c_w_148;
wire [1505:0] c_w_149;
wire [1505:0] c_w_150;
wire [1505:0] c_w_151;
wire [1505:0] c_w_152;
wire [1505:0] c_w_153;
wire [1505:0] c_w_154;
wire [1505:0] c_w_155;
wire [1505:0] c_w_156;
wire [1505:0] c_w_157;
wire [1505:0] c_w_158;
wire [1505:0] c_w_159;
wire [1505:0] c_w_160;
wire [1505:0] c_w_161;
wire [1505:0] c_w_162;
wire [1505:0] c_w_163;
wire [1505:0] c_w_164;
wire [1505:0] c_w_165;
wire [1505:0] c_w_166;
wire [1505:0] c_w_167;
wire [1505:0] c_w_168;
wire [1505:0] c_w_169;
wire [1505:0] c_w_170;
wire [1505:0] c_w_171;
wire [1505:0] c_w_172;
wire [1505:0] c_w_173;
wire [1505:0] c_w_174;
wire [1505:0] c_w_175;
wire [1505:0] c_w_176;
wire [1505:0] c_w_177;
wire [1505:0] c_w_178;
wire [1505:0] c_w_179;
wire [1505:0] c_w_180;
wire [1505:0] c_w_181;
wire [1505:0] c_w_182;
wire [1505:0] c_w_183;
wire [1505:0] c_w_184;
wire [1505:0] c_w_185;
wire [1505:0] c_w_186;
wire [1505:0] c_w_187;
wire [1505:0] c_w_188;
wire [1505:0] c_w_189;
wire [1505:0] c_w_190;
wire [1505:0] c_w_191;
wire [1505:0] c_w_192;
wire [1505:0] c_w_193;
wire [1505:0] c_w_194;
wire [1505:0] c_w_195;
wire [1505:0] c_w_196;
wire [1505:0] c_w_197;
wire [1505:0] c_w_198;
wire [1505:0] c_w_199;
wire [1505:0] c_w_200;
wire [1505:0] c_w_201;
wire [1505:0] c_w_202;
wire [1505:0] c_w_203;
wire [1505:0] c_w_204;
wire [1505:0] c_w_205;
wire [1505:0] c_w_206;
wire [1505:0] c_w_207;
wire [1505:0] c_w_208;
wire [1505:0] c_w_209;
wire [1505:0] c_w_210;
wire [1505:0] c_w_211;
wire [1505:0] c_w_212;
wire [1505:0] c_w_213;
wire [1505:0] c_w_214;
wire [1505:0] c_w_215;
wire [1505:0] c_w_216;
wire [1505:0] c_w_217;
wire [1505:0] c_w_218;
wire [1505:0] c_w_219;
wire [1505:0] c_w_220;
wire [1505:0] c_w_221;
wire [1505:0] c_w_222;
wire [1505:0] c_w_223;
wire [1505:0] c_w_224;
wire [1505:0] c_w_225;
wire [1505:0] c_w_226;
wire [1505:0] c_w_227;
wire [1505:0] c_w_228;
wire [1505:0] c_w_229;
wire [1505:0] c_w_230;
wire [1505:0] c_w_231;
wire [1505:0] c_w_232;
wire [1505:0] c_w_233;
wire [1505:0] c_w_234;
wire [1505:0] c_w_235;
wire [1505:0] c_w_236;
wire [1505:0] c_w_237;
wire [1505:0] c_w_238;
wire [1505:0] c_w_239;
wire [1505:0] c_w_240;
wire [1505:0] c_w_241;
wire [1505:0] c_w_242;
wire [1505:0] c_w_243;
wire [1505:0] c_w_244;
wire [1505:0] c_w_245;
wire [1505:0] c_w_246;
wire [1505:0] c_w_247;
wire [1505:0] c_w_248;
wire [1505:0] c_w_249;
wire [1505:0] c_w_250;
wire [1505:0] c_w_251;
wire [1505:0] c_w_252;
wire [1505:0] c_w_253;
wire [1505:0] c_w_254;
wire [1505:0] c_w_255;
wire [1505:0] c_w_256;
wire [1505:0] c_w_257;
wire [1505:0] c_w_258;
wire [1505:0] c_w_259;
wire [1505:0] c_w_260;
wire [1505:0] c_w_261;
wire [1505:0] c_w_262;
wire [1505:0] c_w_263;
wire [1505:0] c_w_264;
wire [1505:0] c_w_265;
wire [1505:0] c_w_266;
wire [1505:0] c_w_267;
wire [1505:0] c_w_268;
wire [1505:0] c_w_269;
wire [1505:0] c_w_270;
wire [1505:0] c_w_271;
wire [1505:0] c_w_272;
wire [1505:0] c_w_273;
wire [1505:0] c_w_274;
wire [1505:0] c_w_275;
wire [1505:0] c_w_276;
wire [1505:0] c_w_277;
wire [1505:0] c_w_278;
wire [1505:0] c_w_279;
wire [1505:0] c_w_280;
wire [1505:0] c_w_281;
wire [1505:0] c_w_282;
wire [1505:0] c_w_283;
wire [1505:0] c_w_284;
wire [1505:0] c_w_285;
wire [1505:0] c_w_286;
wire [1505:0] c_w_287;
wire [1505:0] c_w_288;
wire [1505:0] c_w_289;
wire [1505:0] c_w_290;
wire [1505:0] c_w_291;
wire [1505:0] c_w_292;
wire [1505:0] c_w_293;
wire [1505:0] c_w_294;
wire [1505:0] c_w_295;
wire [1505:0] c_w_296;
wire [1505:0] c_w_297;
wire [1505:0] c_w_298;
wire [1505:0] c_w_299;
wire [1505:0] c_w_300;
wire [1505:0] c_w_301;
wire [1505:0] c_w_302;
wire [1505:0] c_w_303;
wire [1505:0] c_w_304;
wire [1505:0] c_w_305;
wire [1505:0] c_w_306;
wire [1505:0] c_w_307;
wire [1505:0] c_w_308;
wire [1505:0] c_w_309;
wire [1505:0] c_w_310;
wire [1505:0] c_w_311;
wire [1505:0] c_w_312;
wire [1505:0] c_w_313;
wire [1505:0] c_w_314;
wire [1505:0] c_w_315;
wire [1505:0] c_w_316;
wire [1505:0] c_w_317;
wire [1505:0] c_w_318;
wire [1505:0] c_w_319;
wire [1505:0] c_w_320;
wire [1505:0] c_w_321;
wire [1505:0] c_w_322;
wire [1505:0] c_w_323;
wire [1505:0] c_w_324;
wire [1505:0] c_w_325;
wire [1505:0] c_w_326;
wire [1505:0] c_w_327;
wire [1505:0] c_w_328;
wire [1505:0] c_w_329;
wire [1505:0] c_w_330;
wire [1505:0] c_w_331;
wire [1505:0] c_w_332;
wire [1505:0] c_w_333;
wire [1505:0] c_w_334;
wire [1505:0] c_w_335;
wire [1505:0] c_w_336;
wire [1505:0] c_w_337;
wire [1505:0] c_w_338;
wire [1505:0] c_w_339;
wire [1505:0] c_w_340;
wire [1505:0] c_w_341;
wire [1505:0] c_w_342;
wire [1505:0] c_w_343;
wire [1505:0] c_w_344;
wire [1505:0] c_w_345;
wire [1505:0] c_w_346;
wire [1505:0] c_w_347;
wire [1505:0] c_w_348;
wire [1505:0] c_w_349;
wire [1505:0] c_w_350;
wire [1505:0] c_w_351;
wire [1505:0] c_w_352;
wire [1505:0] c_w_353;
wire [1505:0] c_w_354;
wire [1505:0] c_w_355;
wire [1505:0] c_w_356;
wire [1505:0] c_w_357;
wire [1505:0] c_w_358;
wire [1505:0] c_w_359;
wire [1505:0] c_w_360;
wire [1505:0] c_w_361;
wire [1505:0] c_w_362;
wire [1505:0] c_w_363;
wire [1505:0] c_w_364;
wire [1505:0] c_w_365;
wire [1505:0] c_w_366;
wire [1505:0] c_w_367;
wire [1505:0] c_w_368;
wire [1505:0] c_w_369;
wire [1505:0] c_w_370;
wire [1505:0] c_w_371;
wire [1505:0] c_w_372;
wire [1505:0] c_w_373;
wire [1505:0] c_w_374;
wire [1505:0] c_w_375;
wire [1505:0] c_w_376;
wire [1505:0] c_w_377;
wire [1505:0] c_w_378;
wire [1505:0] c_w_379;
wire [1505:0] c_w_380;
wire [1505:0] c_w_381;
wire [1505:0] c_w_382;
wire [1505:0] c_w_383;
wire [1505:0] c_w_384;
wire [1505:0] c_w_385;
wire [1505:0] c_w_386;
wire [1505:0] c_w_387;
wire [1505:0] c_w_388;
wire [1505:0] c_w_389;
wire [1505:0] c_w_390;
wire [1505:0] c_w_391;
wire [1505:0] c_w_392;
wire [1505:0] c_w_393;
wire [1505:0] c_w_394;
wire [1505:0] c_w_395;
wire [1505:0] c_w_396;
wire [1505:0] c_w_397;
wire [1505:0] c_w_398;
wire [1505:0] c_w_399;
wire [1505:0] c_w_400;
wire [1505:0] c_w_401;
wire [1505:0] c_w_402;
wire [1505:0] c_w_403;
wire [1505:0] c_w_404;
wire [1505:0] c_w_405;
wire [1505:0] c_w_406;
wire [1505:0] c_w_407;
wire [1505:0] c_w_408;
wire [1505:0] c_w_409;
wire [1505:0] c_w_410;
wire [1505:0] c_w_411;
wire [1505:0] c_w_412;
wire [1505:0] c_w_413;
wire [1505:0] c_w_414;
wire [1505:0] c_w_415;
wire [1505:0] c_w_416;
wire [1505:0] c_w_417;
wire [1505:0] c_w_418;
wire [1505:0] c_w_419;
wire [1505:0] c_w_420;
wire [1505:0] c_w_421;
wire [1505:0] c_w_422;
wire [1505:0] c_w_423;
wire [1505:0] c_w_424;
wire [1505:0] c_w_425;
wire [1505:0] c_w_426;
wire [1505:0] c_w_427;
wire [1505:0] c_w_428;
wire [1505:0] c_w_429;
wire [1505:0] c_w_430;
wire [1505:0] c_w_431;
wire [1505:0] c_w_432;
wire [1505:0] c_w_433;
wire [1505:0] c_w_434;
wire [1505:0] c_w_435;
wire [1505:0] c_w_436;
wire [1505:0] c_w_437;
wire [1505:0] c_w_438;
wire [1505:0] c_w_439;
wire [1505:0] c_w_440;
wire [1505:0] c_w_441;
wire [1505:0] c_w_442;
wire [1505:0] c_w_443;
wire [1505:0] c_w_444;
wire [1505:0] c_w_445;
wire [1505:0] c_w_446;
wire [1505:0] c_w_447;
wire [1505:0] c_w_448;
wire [1505:0] c_w_449;
wire [1505:0] c_w_450;
wire [1505:0] c_w_451;
wire [1505:0] c_w_452;
wire [1505:0] c_w_453;
wire [1505:0] c_w_454;
wire [1505:0] c_w_455;
wire [1505:0] c_w_456;
wire [1505:0] c_w_457;
wire [1505:0] c_w_458;
wire [1505:0] c_w_459;
wire [1505:0] c_w_460;
wire [1505:0] c_w_461;
wire [1505:0] c_w_462;
wire [1505:0] c_w_463;
wire [1505:0] c_w_464;
wire [1505:0] c_w_465;
wire [1505:0] c_w_466;
wire [1505:0] c_w_467;
wire [1505:0] c_w_468;
wire [1505:0] c_w_469;
wire [1505:0] c_w_470;
wire [1505:0] c_w_471;
wire [1505:0] c_w_472;
wire [1505:0] c_w_473;
wire [1505:0] c_w_474;
wire [1505:0] c_w_475;
wire [1505:0] c_w_476;
wire [1505:0] c_w_477;
wire [1505:0] c_w_478;
wire [1505:0] c_w_479;
wire [1505:0] c_w_480;
wire [1505:0] c_w_481;
wire [1505:0] c_w_482;
wire [1505:0] c_w_483;
wire [1505:0] c_w_484;
wire [1505:0] c_w_485;
wire [1505:0] c_w_486;
wire [1505:0] c_w_487;
wire [1505:0] c_w_488;
wire [1505:0] c_w_489;
wire [1505:0] c_w_490;
wire [1505:0] c_w_491;
wire [1505:0] c_w_492;
wire [1505:0] c_w_493;
wire [1505:0] c_w_494;
wire [1505:0] c_w_495;
wire [1505:0] c_w_496;
wire [1505:0] c_w_497;
wire [1505:0] c_w_498;
wire [1505:0] c_w_499;
wire [1505:0] c_w_500;
wire [1505:0] c_w_501;
wire [1505:0] c_w_502;
wire [1505:0] c_w_503;
wire [1505:0] c_w_504;
wire [1505:0] c_w_505;
wire [1505:0] c_w_506;
wire [1505:0] c_w_507;
wire [1505:0] c_w_508;
wire [1505:0] c_w_509;
wire [1505:0] c_w_510;
wire [1505:0] c_w_511;
wire [1505:0] c_w_512;
wire [1505:0] c_w_513;
wire [1505:0] c_w_514;
wire [1505:0] c_w_515;
wire [1505:0] c_w_516;
wire [1505:0] c_w_517;
wire [1505:0] c_w_518;
wire [1505:0] c_w_519;
wire [1505:0] c_w_520;
wire [1505:0] c_w_521;
wire [1505:0] c_w_522;
wire [1505:0] c_w_523;
wire [1505:0] c_w_524;
wire [1505:0] c_w_525;
wire [1505:0] c_w_526;
wire [1505:0] c_w_527;
wire [1505:0] c_w_528;
wire [1505:0] c_w_529;
wire [1505:0] c_w_530;
wire [1505:0] c_w_531;
wire [1505:0] c_w_532;
wire [1505:0] c_w_533;
wire [1505:0] c_w_534;
wire [1505:0] c_w_535;
wire [1505:0] c_w_536;
wire [1505:0] c_w_537;
wire [1505:0] c_w_538;
wire [1505:0] c_w_539;
wire [1505:0] c_w_540;
wire [1505:0] c_w_541;
wire [1505:0] c_w_542;
wire [1505:0] c_w_543;
wire [1505:0] c_w_544;
wire [1505:0] c_w_545;
wire [1505:0] c_w_546;
wire [1505:0] c_w_547;
wire [1505:0] c_w_548;
wire [1505:0] c_w_549;
wire [1505:0] c_w_550;
wire [1505:0] c_w_551;
wire [1505:0] c_w_552;
wire [1505:0] c_w_553;
wire [1505:0] c_w_554;
wire [1505:0] c_w_555;
wire [1505:0] c_w_556;
wire [1505:0] c_w_557;
wire [1505:0] c_w_558;
wire [1505:0] c_w_559;
wire [1505:0] c_w_560;
wire [1505:0] c_w_561;
wire [1505:0] c_w_562;
wire [1505:0] c_w_563;
wire [1505:0] c_w_564;
wire [1505:0] c_w_565;
wire [1505:0] c_w_566;
wire [1505:0] c_w_567;
wire [1505:0] c_w_568;
wire [1505:0] c_w_569;
wire [1505:0] c_w_570;
wire [1505:0] c_w_571;
wire [1505:0] c_w_572;
wire [1505:0] c_w_573;
wire [1505:0] c_w_574;
wire [1505:0] c_w_575;
wire [1505:0] c_w_576;
wire [1505:0] c_w_577;
wire [1505:0] c_w_578;
wire [1505:0] c_w_579;
wire [1505:0] c_w_580;
wire [1505:0] c_w_581;
wire [1505:0] c_w_582;
wire [1505:0] c_w_583;
wire [1505:0] c_w_584;
wire [1505:0] c_w_585;
wire [1505:0] c_w_586;
wire [1505:0] c_w_587;
wire [1505:0] c_w_588;
wire [1505:0] c_w_589;
wire [1505:0] c_w_590;
wire [1505:0] c_w_591;
wire [1505:0] c_w_592;
wire [1505:0] c_w_593;
wire [1505:0] c_w_594;
wire [1505:0] c_w_595;
wire [1505:0] c_w_596;
wire [1505:0] c_w_597;
wire [1505:0] c_w_598;
wire [1505:0] c_w_599;
wire [1505:0] c_w_600;
wire [1505:0] c_w_601;
wire [1505:0] c_w_602;
wire [1505:0] c_w_603;
wire [1505:0] c_w_604;
wire [1505:0] c_w_605;
wire [1505:0] c_w_606;
wire [1505:0] c_w_607;
wire [1505:0] c_w_608;
wire [1505:0] c_w_609;
wire [1505:0] c_w_610;
wire [1505:0] c_w_611;
wire [1505:0] c_w_612;
wire [1505:0] c_w_613;
wire [1505:0] c_w_614;
wire [1505:0] c_w_615;
wire [1505:0] c_w_616;
wire [1505:0] c_w_617;
wire [1505:0] c_w_618;
wire [1505:0] c_w_619;
wire [1505:0] c_w_620;
wire [1505:0] c_w_621;
wire [1505:0] c_w_622;
wire [1505:0] c_w_623;
wire [1505:0] c_w_624;
wire [1505:0] c_w_625;
wire [1505:0] c_w_626;
wire [1505:0] c_w_627;
wire [1505:0] c_w_628;
wire [1505:0] c_w_629;
wire [1505:0] c_w_630;
wire [1505:0] c_w_631;
wire [1505:0] c_w_632;
wire [1505:0] c_w_633;
wire [1505:0] c_w_634;
wire [1505:0] c_w_635;
wire [1505:0] c_w_636;
wire [1505:0] c_w_637;
wire [1505:0] c_w_638;
wire [1505:0] c_w_639;
wire [1505:0] c_w_640;
wire [1505:0] c_w_641;
wire [1505:0] c_w_642;
wire [1505:0] c_w_643;
wire [1505:0] c_w_644;
wire [1505:0] c_w_645;
wire [1505:0] c_w_646;
wire [1505:0] c_w_647;
wire [1505:0] c_w_648;
wire [1505:0] c_w_649;
wire [1505:0] c_w_650;
wire [1505:0] c_w_651;
wire [1505:0] c_w_652;
wire [1505:0] c_w_653;
wire [1505:0] c_w_654;
wire [1505:0] c_w_655;
wire [1505:0] c_w_656;
wire [1505:0] c_w_657;
wire [1505:0] c_w_658;
wire [1505:0] c_w_659;
wire [1505:0] c_w_660;
wire [1505:0] c_w_661;
wire [1505:0] c_w_662;
wire [1505:0] c_w_663;
wire [1505:0] c_w_664;
wire [1505:0] c_w_665;
wire [1505:0] c_w_666;
wire [1505:0] c_w_667;
wire [1505:0] c_w_668;
wire [1505:0] c_w_669;
wire [1505:0] c_w_670;
wire [1505:0] c_w_671;
wire [1505:0] c_w_672;
wire [1505:0] c_w_673;
wire [1505:0] c_w_674;
wire [1505:0] c_w_675;
wire [1505:0] c_w_676;
wire [1505:0] c_w_677;
wire [1505:0] c_w_678;
wire [1505:0] c_w_679;
wire [1505:0] c_w_680;
wire [1505:0] c_w_681;
wire [1505:0] c_w_682;
wire [1505:0] c_w_683;
wire [1505:0] c_w_684;
wire [1505:0] c_w_685;
wire [1505:0] c_w_686;
wire [1505:0] c_w_687;
wire [1505:0] c_w_688;
wire [1505:0] c_w_689;
wire [1505:0] c_w_690;
wire [1505:0] c_w_691;
wire [1505:0] c_w_692;
wire [1505:0] c_w_693;
wire [1505:0] c_w_694;
wire [1505:0] c_w_695;
wire [1505:0] c_w_696;
wire [1505:0] c_w_697;
wire [1505:0] c_w_698;
wire [1505:0] c_w_699;
wire [1505:0] c_w_700;
wire [1505:0] c_w_701;
wire [1505:0] c_w_702;
wire [1505:0] c_w_703;
wire [1505:0] c_w_704;
wire [1505:0] c_w_705;
wire [1505:0] c_w_706;
wire [1505:0] c_w_707;
wire [1505:0] c_w_708;
wire [1505:0] c_w_709;
wire [1505:0] c_w_710;
wire [1505:0] c_w_711;
wire [1505:0] c_w_712;
wire [1505:0] c_w_713;
wire [1505:0] c_w_714;
wire [1505:0] c_w_715;
wire [1505:0] c_w_716;
wire [1505:0] c_w_717;
wire [1505:0] c_w_718;
wire [1505:0] c_w_719;
wire [1505:0] c_w_720;
wire [1505:0] c_w_721;
wire [1505:0] c_w_722;
wire [1505:0] c_w_723;
wire [1505:0] c_w_724;
wire [1505:0] c_w_725;
wire [1505:0] c_w_726;
wire [1505:0] c_w_727;
wire [1505:0] c_w_728;
wire [1505:0] c_w_729;
wire [1505:0] c_w_730;
wire [1505:0] c_w_731;
wire [1505:0] c_w_732;
wire [1505:0] c_w_733;
wire [1505:0] c_w_734;
wire [1505:0] c_w_735;
wire [1505:0] c_w_736;
wire [1505:0] c_w_737;
wire [1505:0] c_w_738;
wire [1505:0] c_w_739;
wire [1505:0] c_w_740;
wire [1505:0] c_w_741;
wire [1505:0] c_w_742;
wire [1505:0] c_w_743;
wire [1505:0] c_w_744;
wire [1505:0] c_w_745;
wire [1505:0] c_w_746;
wire [1505:0] c_w_747;
wire [1505:0] c_w_748;
wire [1505:0] c_w_749;
wire [1505:0] c_w_750;
wire [1505:0] c_w_751;
wire [1505:0] c_w_752;
wire [1505:0] c_w_753;
wire [1505:0] c_w_754;
wire [1505:0] c_w_755;
wire [1505:0] c_w_756;
wire [1505:0] c_w_757;
wire [1505:0] c_w_758;
wire [1505:0] c_w_759;
wire [1505:0] c_w_760;
wire [1505:0] c_w_761;
wire [1505:0] c_w_762;
wire [1505:0] c_w_763;
wire [1505:0] c_w_764;
wire [1505:0] c_w_765;
wire [1505:0] c_w_766;
wire [1505:0] c_w_767;
wire [1505:0] c_w_768;
wire [1505:0] c_w_769;
wire [1505:0] c_w_770;
wire [1505:0] c_w_771;
wire [1505:0] c_w_772;
wire [1505:0] c_w_773;
wire [1505:0] c_w_774;
wire [1505:0] c_w_775;
wire [1505:0] c_w_776;
wire [1505:0] c_w_777;
wire [1505:0] c_w_778;
wire [1505:0] c_w_779;
wire [1505:0] c_w_780;
wire [1505:0] c_w_781;
wire [1505:0] c_w_782;
wire [1505:0] c_w_783;
wire [1505:0] c_w_784;
wire [1505:0] c_w_785;
wire [1505:0] c_w_786;
wire [1505:0] c_w_787;
wire [1505:0] c_w_788;
wire [1505:0] c_w_789;
wire [1505:0] c_w_790;
wire [1505:0] c_w_791;
wire [1505:0] c_w_792;
wire [1505:0] c_w_793;
wire [1505:0] c_w_794;
wire [1505:0] c_w_795;
wire [1505:0] c_w_796;
wire [1505:0] c_w_797;
wire [1505:0] c_w_798;
wire [1505:0] c_w_799;
wire [1505:0] c_w_800;
wire [1505:0] c_w_801;
wire [1505:0] c_w_802;
wire [1505:0] c_w_803;
wire [1505:0] c_w_804;
wire [1505:0] c_w_805;
wire [1505:0] c_w_806;
wire [1505:0] c_w_807;
wire [1505:0] c_w_808;
wire [1505:0] c_w_809;
wire [1505:0] c_w_810;
wire [1505:0] c_w_811;
wire [1505:0] c_w_812;
wire [1505:0] c_w_813;
wire [1505:0] c_w_814;
wire [1505:0] c_w_815;
wire [1505:0] c_w_816;
wire [1505:0] c_w_817;
wire [1505:0] c_w_818;
wire [1505:0] c_w_819;
wire [1505:0] c_w_820;
wire [1505:0] c_w_821;
wire [1505:0] c_w_822;
wire [1505:0] c_w_823;
wire [1505:0] c_w_824;
wire [1505:0] c_w_825;
wire [1505:0] c_w_826;
wire [1505:0] c_w_827;
wire [1505:0] c_w_828;
wire [1505:0] c_w_829;
wire [1505:0] c_w_830;
wire [1505:0] c_w_831;
wire [1505:0] c_w_832;
wire [1505:0] c_w_833;
wire [1505:0] c_w_834;
wire [1505:0] c_w_835;
wire [1505:0] c_w_836;
wire [1505:0] c_w_837;
wire [1505:0] c_w_838;
wire [1505:0] c_w_839;
wire [1505:0] c_w_840;
wire [1505:0] c_w_841;
wire [1505:0] c_w_842;
wire [1505:0] c_w_843;
wire [1505:0] c_w_844;
wire [1505:0] c_w_845;
wire [1505:0] c_w_846;
wire [1505:0] c_w_847;
wire [1505:0] c_w_848;
wire [1505:0] c_w_849;
wire [1505:0] c_w_850;
wire [1505:0] c_w_851;
wire [1505:0] c_w_852;
wire [1505:0] c_w_853;
wire [1505:0] c_w_854;
wire [1505:0] c_w_855;
wire [1505:0] c_w_856;
wire [1505:0] c_w_857;
wire [1505:0] c_w_858;
wire [1505:0] c_w_859;
wire [1505:0] c_w_860;
wire [1505:0] c_w_861;
wire [1505:0] c_w_862;
wire [1505:0] c_w_863;
wire [1505:0] c_w_864;
wire [1505:0] c_w_865;
wire [1505:0] c_w_866;
wire [1505:0] c_w_867;
wire [1505:0] c_w_868;
wire [1505:0] c_w_869;
wire [1505:0] c_w_870;
wire [1505:0] c_w_871;
wire [1505:0] c_w_872;
wire [1505:0] c_w_873;
wire [1505:0] c_w_874;
wire [1505:0] c_w_875;
wire [1505:0] c_w_876;
wire [1505:0] c_w_877;
wire [1505:0] c_w_878;
wire [1505:0] c_w_879;
wire [1505:0] c_w_880;
wire [1505:0] c_w_881;
wire [1505:0] c_w_882;
wire [1505:0] c_w_883;
wire [1505:0] c_w_884;
wire [1505:0] c_w_885;
wire [1505:0] c_w_886;
wire [1505:0] c_w_887;
wire [1505:0] c_w_888;
wire [1505:0] c_w_889;
wire [1505:0] c_w_890;
wire [1505:0] c_w_891;
wire [1505:0] c_w_892;
wire [1505:0] c_w_893;
wire [1505:0] c_w_894;
wire [1505:0] c_w_895;
wire [1505:0] c_w_896;
wire [1505:0] c_w_897;
wire [1505:0] c_w_898;
wire [1505:0] c_w_899;
wire [1505:0] c_w_900;
wire [1505:0] c_w_901;
wire [1505:0] c_w_902;
wire [1505:0] c_w_903;
wire [1505:0] c_w_904;
wire [1505:0] c_w_905;
wire [1505:0] c_w_906;
wire [1505:0] c_w_907;
wire [1505:0] c_w_908;
wire [1505:0] c_w_909;
wire [1505:0] c_w_910;
wire [1505:0] c_w_911;
wire [1505:0] c_w_912;
wire [1505:0] c_w_913;
wire [1505:0] c_w_914;
wire [1505:0] c_w_915;
wire [1505:0] c_w_916;
wire [1505:0] c_w_917;
wire [1505:0] c_w_918;
wire [1505:0] c_w_919;
wire [1505:0] c_w_920;
wire [1505:0] c_w_921;
wire [1505:0] c_w_922;
wire [1505:0] c_w_923;
wire [1505:0] c_w_924;
wire [1505:0] c_w_925;
wire [1505:0] c_w_926;
wire [1505:0] c_w_927;
wire [1505:0] c_w_928;
wire [1505:0] c_w_929;
wire [1505:0] c_w_930;
wire [1505:0] c_w_931;
wire [1505:0] c_w_932;
wire [1505:0] c_w_933;
wire [1505:0] c_w_934;
wire [1505:0] c_w_935;
wire [1505:0] c_w_936;
wire [1505:0] c_w_937;
wire [1505:0] c_w_938;
wire [1505:0] c_w_939;
wire [1505:0] c_w_940;
wire [1505:0] c_w_941;
wire [1505:0] c_w_942;
wire [1505:0] c_w_943;
wire [1505:0] c_w_944;
wire [1505:0] c_w_945;
wire [1505:0] c_w_946;
wire [1505:0] c_w_947;
wire [1505:0] c_w_948;
wire [1505:0] c_w_949;
wire [1505:0] c_w_950;
wire [1505:0] c_w_951;
wire [1505:0] c_w_952;
wire [1505:0] c_w_953;
wire [1505:0] c_w_954;
wire [1505:0] c_w_955;
wire [1505:0] c_w_956;
wire [1505:0] c_w_957;
wire [1505:0] c_w_958;
wire [1505:0] c_w_959;
wire [1505:0] c_w_960;
wire [1505:0] c_w_961;
wire [1505:0] c_w_962;
wire [1505:0] c_w_963;
wire [1505:0] c_w_964;
wire [1505:0] c_w_965;
wire [1505:0] c_w_966;
wire [1505:0] c_w_967;
wire [1505:0] c_w_968;
wire [1505:0] c_w_969;
wire [1505:0] c_w_970;
wire [1505:0] c_w_971;
wire [1505:0] c_w_972;
wire [1505:0] c_w_973;
wire [1505:0] c_w_974;
wire [1505:0] c_w_975;
wire [1505:0] c_w_976;
wire [1505:0] c_w_977;
wire [1505:0] c_w_978;
wire [1505:0] c_w_979;
wire [1505:0] c_w_980;
wire [1505:0] c_w_981;
wire [1505:0] c_w_982;
wire [1505:0] c_w_983;
wire [1505:0] c_w_984;
wire [1505:0] c_w_985;
wire [1505:0] c_w_986;
wire [1505:0] c_w_987;
wire [1505:0] c_w_988;
wire [1505:0] c_w_989;
wire [1505:0] c_w_990;
wire [1505:0] c_w_991;
wire [1505:0] c_w_992;
wire [1505:0] c_w_993;
wire [1505:0] c_w_994;
wire [1505:0] c_w_995;
wire [1505:0] c_w_996;
wire [1505:0] c_w_997;
wire [1505:0] c_w_998;
wire [1505:0] c_w_999;
wire [1505:0] c_w_1000;
wire [1505:0] c_w_1001;
wire [1505:0] c_w_1002;
wire [1505:0] c_w_1003;
wire [1505:0] c_w_1004;
wire [1505:0] c_w_1005;
wire [1505:0] c_w_1006;
wire [1505:0] c_w_1007;
wire [1505:0] c_w_1008;
wire [1505:0] c_w_1009;
wire [1505:0] c_w_1010;
wire [1505:0] c_w_1011;
wire [1505:0] c_w_1012;
wire [1505:0] c_w_1013;
wire [1505:0] c_w_1014;
wire [1505:0] c_w_1015;
wire [1505:0] c_w_1016;
wire [1505:0] c_w_1017;
wire [1505:0] c_w_1018;
wire [1505:0] c_w_1019;
wire [1505:0] c_w_1020;
wire [1505:0] c_w_1021;
wire [1505:0] c_w_1022;
wire [1505:0] c_w_1023;
wire [1505:0] c_w_1024;
wire [1505:0] c_w_1025;
wire [1505:0] c_w_1026;
wire [1505:0] c_w_1027;
wire [1505:0] c_w_1028;
wire [1505:0] c_w_1029;
wire [1505:0] c_w_1030;
wire [1505:0] c_w_1031;
wire [1505:0] c_w_1032;
wire [1505:0] c_w_1033;
wire [1505:0] c_w_1034;
wire [1505:0] c_w_1035;
wire [1505:0] c_w_1036;
wire [1505:0] c_w_1037;
wire [1505:0] c_w_1038;
wire [1505:0] c_w_1039;
wire [1505:0] c_w_1040;
wire [1505:0] c_w_1041;
wire [1505:0] c_w_1042;
wire [1505:0] c_w_1043;
wire [1505:0] c_w_1044;
wire [1505:0] c_w_1045;
wire [1505:0] c_w_1046;
wire [1505:0] c_w_1047;
wire [1505:0] c_w_1048;
wire [1505:0] c_w_1049;
wire [1505:0] c_w_1050;
wire [1505:0] c_w_1051;
wire [1505:0] c_w_1052;
wire [1505:0] c_w_1053;
wire [1505:0] c_w_1054;
wire [1505:0] c_w_1055;
wire [1505:0] c_w_1056;
wire [1505:0] c_w_1057;
wire [1505:0] c_w_1058;
wire [1505:0] c_w_1059;
wire [1505:0] c_w_1060;
wire [1505:0] c_w_1061;
wire [1505:0] c_w_1062;
wire [1505:0] c_w_1063;
wire [1505:0] c_w_1064;
wire [1505:0] c_w_1065;
wire [1505:0] c_w_1066;
wire [1505:0] c_w_1067;
wire [1505:0] c_w_1068;
wire [1505:0] c_w_1069;
wire [1505:0] c_w_1070;
wire [1505:0] c_w_1071;
wire [1505:0] c_w_1072;
wire [1505:0] c_w_1073;
wire [1505:0] c_w_1074;
wire [1505:0] c_w_1075;
wire [1505:0] c_w_1076;
wire [1505:0] c_w_1077;
wire [1505:0] c_w_1078;
wire [1505:0] c_w_1079;
wire [1505:0] c_w_1080;
wire [1505:0] c_w_1081;
wire [1505:0] c_w_1082;
wire [1505:0] c_w_1083;
wire [1505:0] c_w_1084;
wire [1505:0] c_w_1085;
wire [1505:0] c_w_1086;
wire [1505:0] c_w_1087;
wire [1505:0] c_w_1088;
wire [1505:0] c_w_1089;
wire [1505:0] c_w_1090;
wire [1505:0] c_w_1091;
wire [1505:0] c_w_1092;
wire [1505:0] c_w_1093;
wire [1505:0] c_w_1094;
wire [1505:0] c_w_1095;
wire [1505:0] c_w_1096;
wire [1505:0] c_w_1097;
wire [1505:0] c_w_1098;
wire [1505:0] c_w_1099;
wire [1505:0] c_w_1100;
wire [1505:0] c_w_1101;
wire [1505:0] c_w_1102;
wire [1505:0] c_w_1103;
wire [1505:0] c_w_1104;
wire [1505:0] c_w_1105;
wire [1505:0] c_w_1106;
wire [1505:0] c_w_1107;
wire [1505:0] c_w_1108;
wire [1505:0] c_w_1109;
wire [1505:0] c_w_1110;
wire [1505:0] c_w_1111;
wire [1505:0] c_w_1112;
wire [1505:0] c_w_1113;
wire [1505:0] c_w_1114;
wire [1505:0] c_w_1115;
wire [1505:0] c_w_1116;
wire [1505:0] c_w_1117;
wire [1505:0] c_w_1118;
wire [1505:0] c_w_1119;
wire [1505:0] c_w_1120;
wire [1505:0] c_w_1121;
wire [1505:0] c_w_1122;
wire [1505:0] c_w_1123;
wire [1505:0] c_w_1124;
wire [1505:0] c_w_1125;
wire [1505:0] c_w_1126;
wire [1505:0] c_w_1127;
wire [1505:0] c_w_1128;
wire [1505:0] c_w_1129;
wire [1505:0] c_w_1130;
wire [1505:0] c_w_1131;
wire [1505:0] c_w_1132;
wire [1505:0] c_w_1133;
wire [1505:0] c_w_1134;
wire [1505:0] c_w_1135;
wire [1505:0] c_w_1136;
wire [1505:0] c_w_1137;
wire [1505:0] c_w_1138;
wire [1505:0] c_w_1139;
wire [1505:0] c_w_1140;
wire [1505:0] c_w_1141;
wire [1505:0] c_w_1142;
wire [1505:0] c_w_1143;
wire [1505:0] c_w_1144;
wire [1505:0] c_w_1145;
wire [1505:0] c_w_1146;
wire [1505:0] c_w_1147;
wire [1505:0] c_w_1148;
wire [1505:0] c_w_1149;
wire [1505:0] c_w_1150;
wire [1505:0] c_w_1151;
wire [1505:0] c_w_1152;
wire [1505:0] c_w_1153;
wire [1505:0] c_w_1154;
wire [1505:0] c_w_1155;
wire [1505:0] c_w_1156;
wire [1505:0] c_w_1157;
wire [1505:0] c_w_1158;
wire [1505:0] c_w_1159;
wire [1505:0] c_w_1160;
wire [1505:0] c_w_1161;
wire [1505:0] c_w_1162;
wire [1505:0] c_w_1163;
wire [1505:0] c_w_1164;
wire [1505:0] c_w_1165;
wire [1505:0] c_w_1166;
wire [1505:0] c_w_1167;
wire [1505:0] c_w_1168;
wire [1505:0] c_w_1169;
wire [1505:0] c_w_1170;
wire [1505:0] c_w_1171;
wire [1505:0] c_w_1172;
wire [1505:0] c_w_1173;
wire [1505:0] c_w_1174;
wire [1505:0] c_w_1175;
wire [1505:0] c_w_1176;
wire [1505:0] c_w_1177;
wire [1505:0] c_w_1178;
wire [1505:0] c_w_1179;
wire [1505:0] c_w_1180;
wire [1505:0] c_w_1181;
wire [1505:0] c_w_1182;
wire [1505:0] c_w_1183;
wire [1505:0] c_w_1184;
wire [1505:0] c_w_1185;
wire [1505:0] c_w_1186;
wire [1505:0] c_w_1187;
wire [1505:0] c_w_1188;
wire [1505:0] c_w_1189;
wire [1505:0] c_w_1190;
wire [1505:0] c_w_1191;
wire [1505:0] c_w_1192;
wire [1505:0] c_w_1193;
wire [1505:0] c_w_1194;
wire [1505:0] c_w_1195;
wire [1505:0] c_w_1196;
wire [1505:0] c_w_1197;
wire [1505:0] c_w_1198;
wire [1505:0] c_w_1199;
wire [1505:0] c_w_1200;
wire [1505:0] c_w_1201;
wire [1505:0] c_w_1202;
wire [1505:0] c_w_1203;
wire [1505:0] c_w_1204;
wire [1505:0] c_w_1205;
wire [1505:0] c_w_1206;
wire [1505:0] c_w_1207;
wire [1505:0] c_w_1208;
wire [1505:0] c_w_1209;
wire [1505:0] c_w_1210;
wire [1505:0] c_w_1211;
wire [1505:0] c_w_1212;
wire [1505:0] c_w_1213;
wire [1505:0] c_w_1214;
wire [1505:0] c_w_1215;
wire [1505:0] c_w_1216;
wire [1505:0] c_w_1217;
wire [1505:0] c_w_1218;
wire [1505:0] c_w_1219;
wire [1505:0] c_w_1220;
wire [1505:0] c_w_1221;
wire [1505:0] c_w_1222;
wire [1505:0] c_w_1223;
wire [1505:0] c_w_1224;
wire [1505:0] c_w_1225;
wire [1505:0] c_w_1226;
wire [1505:0] c_w_1227;
wire [1505:0] c_w_1228;
wire [1505:0] c_w_1229;
wire [1505:0] c_w_1230;
wire [1505:0] c_w_1231;
wire [1505:0] c_w_1232;
wire [1505:0] c_w_1233;
wire [1505:0] c_w_1234;
wire [1505:0] c_w_1235;
wire [1505:0] c_w_1236;
wire [1505:0] c_w_1237;
wire [1505:0] c_w_1238;
wire [1505:0] c_w_1239;
wire [1505:0] c_w_1240;
wire [1505:0] c_w_1241;
wire [1505:0] c_w_1242;
wire [1505:0] c_w_1243;
wire [1505:0] c_w_1244;
wire [1505:0] c_w_1245;
wire [1505:0] c_w_1246;
wire [1505:0] c_w_1247;
wire [1505:0] c_w_1248;
wire [1505:0] c_w_1249;
wire [1505:0] c_w_1250;
wire [1505:0] c_w_1251;
wire [1505:0] c_w_1252;
wire [1505:0] c_w_1253;
wire [1505:0] c_w_1254;
wire [1505:0] c_w_1255;
wire [1505:0] c_w_1256;
wire [1505:0] c_w_1257;
wire [1505:0] c_w_1258;
wire [1505:0] c_w_1259;
wire [1505:0] c_w_1260;
wire [1505:0] c_w_1261;
wire [1505:0] c_w_1262;
wire [1505:0] c_w_1263;
wire [1505:0] c_w_1264;
wire [1505:0] c_w_1265;
wire [1505:0] c_w_1266;
wire [1505:0] c_w_1267;
wire [1505:0] c_w_1268;
wire [1505:0] c_w_1269;
wire [1505:0] c_w_1270;
wire [1505:0] c_w_1271;
wire [1505:0] c_w_1272;
wire [1505:0] c_w_1273;
wire [1505:0] c_w_1274;
wire [1505:0] c_w_1275;
wire [1505:0] c_w_1276;
wire [1505:0] c_w_1277;
wire [1505:0] c_w_1278;
wire [1505:0] c_w_1279;
wire [1505:0] c_w_1280;
wire [1505:0] c_w_1281;
wire [1505:0] c_w_1282;
wire [1505:0] c_w_1283;
wire [1505:0] c_w_1284;
wire [1505:0] c_w_1285;
wire [1505:0] c_w_1286;
wire [1505:0] c_w_1287;
wire [1505:0] c_w_1288;
wire [1505:0] c_w_1289;
wire [1505:0] c_w_1290;
wire [1505:0] c_w_1291;
wire [1505:0] c_w_1292;
wire [1505:0] c_w_1293;
wire [1505:0] c_w_1294;
wire [1505:0] c_w_1295;
wire [1505:0] c_w_1296;
wire [1505:0] c_w_1297;
wire [1505:0] c_w_1298;
wire [1505:0] c_w_1299;
wire [1505:0] c_w_1300;
wire [1505:0] c_w_1301;
wire [1505:0] c_w_1302;
wire [1505:0] c_w_1303;
wire [1505:0] c_w_1304;
wire [1505:0] c_w_1305;
wire [1505:0] c_w_1306;
wire [1505:0] c_w_1307;
wire [1505:0] c_w_1308;
wire [1505:0] c_w_1309;
wire [1505:0] c_w_1310;
wire [1505:0] c_w_1311;
wire [1505:0] c_w_1312;
wire [1505:0] c_w_1313;
wire [1505:0] c_w_1314;
wire [1505:0] c_w_1315;
wire [1505:0] c_w_1316;
wire [1505:0] c_w_1317;
wire [1505:0] c_w_1318;
wire [1505:0] c_w_1319;
wire [1505:0] c_w_1320;
wire [1505:0] c_w_1321;
wire [1505:0] c_w_1322;
wire [1505:0] c_w_1323;
wire [1505:0] c_w_1324;
wire [1505:0] c_w_1325;
wire [1505:0] c_w_1326;
wire [1505:0] c_w_1327;
wire [1505:0] c_w_1328;
wire [1505:0] c_w_1329;
wire [1505:0] c_w_1330;
wire [1505:0] c_w_1331;
wire [1505:0] c_w_1332;
wire [1505:0] c_w_1333;
wire [1505:0] c_w_1334;
wire [1505:0] c_w_1335;
wire [1505:0] c_w_1336;
wire [1505:0] c_w_1337;
wire [1505:0] c_w_1338;
wire [1505:0] c_w_1339;
wire [1505:0] c_w_1340;
wire [1505:0] c_w_1341;
wire [1505:0] c_w_1342;
wire [1505:0] c_w_1343;
wire [1505:0] c_w_1344;
wire [1505:0] c_w_1345;
wire [1505:0] c_w_1346;
wire [1505:0] c_w_1347;
wire [1505:0] c_w_1348;
wire [1505:0] c_w_1349;
wire [1505:0] c_w_1350;
wire [1505:0] c_w_1351;
wire [1505:0] c_w_1352;
wire [1505:0] c_w_1353;
wire [1505:0] c_w_1354;
wire [1505:0] c_w_1355;
wire [1505:0] c_w_1356;
wire [1505:0] c_w_1357;
wire [1505:0] c_w_1358;
wire [1505:0] c_w_1359;
wire [1505:0] c_w_1360;
wire [1505:0] c_w_1361;
wire [1505:0] c_w_1362;
wire [1505:0] c_w_1363;
wire [1505:0] c_w_1364;
wire [1505:0] c_w_1365;
wire [1505:0] c_w_1366;
wire [1505:0] c_w_1367;
wire [1505:0] c_w_1368;
wire [1505:0] c_w_1369;
wire [1505:0] c_w_1370;
wire [1505:0] c_w_1371;
wire [1505:0] c_w_1372;
wire [1505:0] c_w_1373;
wire [1505:0] c_w_1374;
wire [1505:0] c_w_1375;
wire [1505:0] c_w_1376;
wire [1505:0] c_w_1377;
wire [1505:0] c_w_1378;
wire [1505:0] c_w_1379;
wire [1505:0] c_w_1380;
wire [1505:0] c_w_1381;
wire [1505:0] c_w_1382;
wire [1505:0] c_w_1383;
wire [1505:0] c_w_1384;
wire [1505:0] c_w_1385;
wire [1505:0] c_w_1386;
wire [1505:0] c_w_1387;
wire [1505:0] c_w_1388;
wire [1505:0] c_w_1389;
wire [1505:0] c_w_1390;
wire [1505:0] c_w_1391;
wire [1505:0] c_w_1392;
wire [1505:0] c_w_1393;
wire [1505:0] c_w_1394;
wire [1505:0] c_w_1395;
wire [1505:0] c_w_1396;
wire [1505:0] c_w_1397;
wire [1505:0] c_w_1398;
wire [1505:0] c_w_1399;
wire [1505:0] c_w_1400;
wire [1505:0] c_w_1401;
wire [1505:0] c_w_1402;
wire [1505:0] c_w_1403;
wire [1505:0] c_w_1404;
wire [1505:0] c_w_1405;
wire [1505:0] c_w_1406;
wire [1505:0] c_w_1407;
wire [1505:0] c_w_1408;
wire [1505:0] c_w_1409;
wire [1505:0] c_w_1410;
wire [1505:0] c_w_1411;
wire [1505:0] c_w_1412;
wire [1505:0] c_w_1413;
wire [1505:0] c_w_1414;
wire [1505:0] c_w_1415;
wire [1505:0] c_w_1416;
wire [1505:0] c_w_1417;
wire [1505:0] c_w_1418;
wire [1505:0] c_w_1419;
wire [1505:0] c_w_1420;
wire [1505:0] c_w_1421;
wire [1505:0] c_w_1422;
wire [1505:0] c_w_1423;
wire [1505:0] c_w_1424;
wire [1505:0] c_w_1425;
wire [1505:0] c_w_1426;
wire [1505:0] c_w_1427;
wire [1505:0] c_w_1428;
wire [1505:0] c_w_1429;
wire [1505:0] c_w_1430;
wire [1505:0] c_w_1431;
wire [1505:0] c_w_1432;
wire [1505:0] c_w_1433;
wire [1505:0] c_w_1434;
wire [1505:0] c_w_1435;
wire [1505:0] c_w_1436;
wire [1505:0] c_w_1437;
wire [1505:0] c_w_1438;
wire [1505:0] c_w_1439;
wire [1505:0] c_w_1440;
wire [1505:0] c_w_1441;
wire [1505:0] c_w_1442;
wire [1505:0] c_w_1443;
wire [1505:0] c_w_1444;
wire [1505:0] c_w_1445;
wire [1505:0] c_w_1446;
wire [1505:0] c_w_1447;
wire [1505:0] c_w_1448;
wire [1505:0] c_w_1449;
wire [1505:0] c_w_1450;
wire [1505:0] c_w_1451;
wire [1505:0] c_w_1452;
wire [1505:0] c_w_1453;
wire [1505:0] c_w_1454;
wire [1505:0] c_w_1455;
wire [1505:0] c_w_1456;
wire [1505:0] c_w_1457;
wire [1505:0] c_w_1458;
wire [1505:0] c_w_1459;
wire [1505:0] c_w_1460;
wire [1505:0] c_w_1461;
wire [1505:0] c_w_1462;
wire [1505:0] c_w_1463;
wire [1505:0] c_w_1464;
wire [1505:0] c_w_1465;
wire [1505:0] c_w_1466;
wire [1505:0] c_w_1467;
wire [1505:0] c_w_1468;
wire [1505:0] c_w_1469;
wire [1505:0] c_w_1470;
wire [1505:0] c_w_1471;
wire [1505:0] c_w_1472;
wire [1505:0] c_w_1473;
wire [1505:0] c_w_1474;
wire [1505:0] c_w_1475;
wire [1505:0] c_w_1476;
wire [1505:0] c_w_1477;
wire [1505:0] c_w_1478;
wire [1505:0] c_w_1479;
wire [1505:0] c_w_1480;
wire [1505:0] c_w_1481;
wire [1505:0] c_w_1482;
wire [1505:0] c_w_1483;
wire [1505:0] c_w_1484;
wire [1505:0] c_w_1485;
wire [1505:0] c_w_1486;
wire [1505:0] c_w_1487;
wire [1505:0] c_w_1488;
wire [1505:0] c_w_1489;
wire [1505:0] c_w_1490;
wire [1505:0] c_w_1491;
wire [1505:0] c_w_1492;
wire [1505:0] c_w_1493;
wire [1505:0] c_w_1494;
wire [1505:0] c_w_1495;
wire [1505:0] c_w_1496;
wire [1505:0] c_w_1497;
wire [1505:0] c_w_1498;
wire [1505:0] c_w_1499;
wire [1505:0] c_w_1500;
wire [1505:0] c_w_1501;
wire [1505:0] c_w_1502;
wire [1505:0] c_w_1503;
wire [1505:0] c_w_1504;
wire [1505:0] c_w_1505;
    
AND_array_1506 AND_array_1506_i0(a,b[0],c_w_0);
AND_array_1506 AND_array_1506_i1(a,b[1],c_w_1);
AND_array_1506 AND_array_1506_i2(a,b[2],c_w_2);
AND_array_1506 AND_array_1506_i3(a,b[3],c_w_3);
AND_array_1506 AND_array_1506_i4(a,b[4],c_w_4);
AND_array_1506 AND_array_1506_i5(a,b[5],c_w_5);
AND_array_1506 AND_array_1506_i6(a,b[6],c_w_6);
AND_array_1506 AND_array_1506_i7(a,b[7],c_w_7);
AND_array_1506 AND_array_1506_i8(a,b[8],c_w_8);
AND_array_1506 AND_array_1506_i9(a,b[9],c_w_9);
AND_array_1506 AND_array_1506_i10(a,b[10],c_w_10);
AND_array_1506 AND_array_1506_i11(a,b[11],c_w_11);
AND_array_1506 AND_array_1506_i12(a,b[12],c_w_12);
AND_array_1506 AND_array_1506_i13(a,b[13],c_w_13);
AND_array_1506 AND_array_1506_i14(a,b[14],c_w_14);
AND_array_1506 AND_array_1506_i15(a,b[15],c_w_15);
AND_array_1506 AND_array_1506_i16(a,b[16],c_w_16);
AND_array_1506 AND_array_1506_i17(a,b[17],c_w_17);
AND_array_1506 AND_array_1506_i18(a,b[18],c_w_18);
AND_array_1506 AND_array_1506_i19(a,b[19],c_w_19);
AND_array_1506 AND_array_1506_i20(a,b[20],c_w_20);
AND_array_1506 AND_array_1506_i21(a,b[21],c_w_21);
AND_array_1506 AND_array_1506_i22(a,b[22],c_w_22);
AND_array_1506 AND_array_1506_i23(a,b[23],c_w_23);
AND_array_1506 AND_array_1506_i24(a,b[24],c_w_24);
AND_array_1506 AND_array_1506_i25(a,b[25],c_w_25);
AND_array_1506 AND_array_1506_i26(a,b[26],c_w_26);
AND_array_1506 AND_array_1506_i27(a,b[27],c_w_27);
AND_array_1506 AND_array_1506_i28(a,b[28],c_w_28);
AND_array_1506 AND_array_1506_i29(a,b[29],c_w_29);
AND_array_1506 AND_array_1506_i30(a,b[30],c_w_30);
AND_array_1506 AND_array_1506_i31(a,b[31],c_w_31);
AND_array_1506 AND_array_1506_i32(a,b[32],c_w_32);
AND_array_1506 AND_array_1506_i33(a,b[33],c_w_33);
AND_array_1506 AND_array_1506_i34(a,b[34],c_w_34);
AND_array_1506 AND_array_1506_i35(a,b[35],c_w_35);
AND_array_1506 AND_array_1506_i36(a,b[36],c_w_36);
AND_array_1506 AND_array_1506_i37(a,b[37],c_w_37);
AND_array_1506 AND_array_1506_i38(a,b[38],c_w_38);
AND_array_1506 AND_array_1506_i39(a,b[39],c_w_39);
AND_array_1506 AND_array_1506_i40(a,b[40],c_w_40);
AND_array_1506 AND_array_1506_i41(a,b[41],c_w_41);
AND_array_1506 AND_array_1506_i42(a,b[42],c_w_42);
AND_array_1506 AND_array_1506_i43(a,b[43],c_w_43);
AND_array_1506 AND_array_1506_i44(a,b[44],c_w_44);
AND_array_1506 AND_array_1506_i45(a,b[45],c_w_45);
AND_array_1506 AND_array_1506_i46(a,b[46],c_w_46);
AND_array_1506 AND_array_1506_i47(a,b[47],c_w_47);
AND_array_1506 AND_array_1506_i48(a,b[48],c_w_48);
AND_array_1506 AND_array_1506_i49(a,b[49],c_w_49);
AND_array_1506 AND_array_1506_i50(a,b[50],c_w_50);
AND_array_1506 AND_array_1506_i51(a,b[51],c_w_51);
AND_array_1506 AND_array_1506_i52(a,b[52],c_w_52);
AND_array_1506 AND_array_1506_i53(a,b[53],c_w_53);
AND_array_1506 AND_array_1506_i54(a,b[54],c_w_54);
AND_array_1506 AND_array_1506_i55(a,b[55],c_w_55);
AND_array_1506 AND_array_1506_i56(a,b[56],c_w_56);
AND_array_1506 AND_array_1506_i57(a,b[57],c_w_57);
AND_array_1506 AND_array_1506_i58(a,b[58],c_w_58);
AND_array_1506 AND_array_1506_i59(a,b[59],c_w_59);
AND_array_1506 AND_array_1506_i60(a,b[60],c_w_60);
AND_array_1506 AND_array_1506_i61(a,b[61],c_w_61);
AND_array_1506 AND_array_1506_i62(a,b[62],c_w_62);
AND_array_1506 AND_array_1506_i63(a,b[63],c_w_63);
AND_array_1506 AND_array_1506_i64(a,b[64],c_w_64);
AND_array_1506 AND_array_1506_i65(a,b[65],c_w_65);
AND_array_1506 AND_array_1506_i66(a,b[66],c_w_66);
AND_array_1506 AND_array_1506_i67(a,b[67],c_w_67);
AND_array_1506 AND_array_1506_i68(a,b[68],c_w_68);
AND_array_1506 AND_array_1506_i69(a,b[69],c_w_69);
AND_array_1506 AND_array_1506_i70(a,b[70],c_w_70);
AND_array_1506 AND_array_1506_i71(a,b[71],c_w_71);
AND_array_1506 AND_array_1506_i72(a,b[72],c_w_72);
AND_array_1506 AND_array_1506_i73(a,b[73],c_w_73);
AND_array_1506 AND_array_1506_i74(a,b[74],c_w_74);
AND_array_1506 AND_array_1506_i75(a,b[75],c_w_75);
AND_array_1506 AND_array_1506_i76(a,b[76],c_w_76);
AND_array_1506 AND_array_1506_i77(a,b[77],c_w_77);
AND_array_1506 AND_array_1506_i78(a,b[78],c_w_78);
AND_array_1506 AND_array_1506_i79(a,b[79],c_w_79);
AND_array_1506 AND_array_1506_i80(a,b[80],c_w_80);
AND_array_1506 AND_array_1506_i81(a,b[81],c_w_81);
AND_array_1506 AND_array_1506_i82(a,b[82],c_w_82);
AND_array_1506 AND_array_1506_i83(a,b[83],c_w_83);
AND_array_1506 AND_array_1506_i84(a,b[84],c_w_84);
AND_array_1506 AND_array_1506_i85(a,b[85],c_w_85);
AND_array_1506 AND_array_1506_i86(a,b[86],c_w_86);
AND_array_1506 AND_array_1506_i87(a,b[87],c_w_87);
AND_array_1506 AND_array_1506_i88(a,b[88],c_w_88);
AND_array_1506 AND_array_1506_i89(a,b[89],c_w_89);
AND_array_1506 AND_array_1506_i90(a,b[90],c_w_90);
AND_array_1506 AND_array_1506_i91(a,b[91],c_w_91);
AND_array_1506 AND_array_1506_i92(a,b[92],c_w_92);
AND_array_1506 AND_array_1506_i93(a,b[93],c_w_93);
AND_array_1506 AND_array_1506_i94(a,b[94],c_w_94);
AND_array_1506 AND_array_1506_i95(a,b[95],c_w_95);
AND_array_1506 AND_array_1506_i96(a,b[96],c_w_96);
AND_array_1506 AND_array_1506_i97(a,b[97],c_w_97);
AND_array_1506 AND_array_1506_i98(a,b[98],c_w_98);
AND_array_1506 AND_array_1506_i99(a,b[99],c_w_99);
AND_array_1506 AND_array_1506_i100(a,b[100],c_w_100);
AND_array_1506 AND_array_1506_i101(a,b[101],c_w_101);
AND_array_1506 AND_array_1506_i102(a,b[102],c_w_102);
AND_array_1506 AND_array_1506_i103(a,b[103],c_w_103);
AND_array_1506 AND_array_1506_i104(a,b[104],c_w_104);
AND_array_1506 AND_array_1506_i105(a,b[105],c_w_105);
AND_array_1506 AND_array_1506_i106(a,b[106],c_w_106);
AND_array_1506 AND_array_1506_i107(a,b[107],c_w_107);
AND_array_1506 AND_array_1506_i108(a,b[108],c_w_108);
AND_array_1506 AND_array_1506_i109(a,b[109],c_w_109);
AND_array_1506 AND_array_1506_i110(a,b[110],c_w_110);
AND_array_1506 AND_array_1506_i111(a,b[111],c_w_111);
AND_array_1506 AND_array_1506_i112(a,b[112],c_w_112);
AND_array_1506 AND_array_1506_i113(a,b[113],c_w_113);
AND_array_1506 AND_array_1506_i114(a,b[114],c_w_114);
AND_array_1506 AND_array_1506_i115(a,b[115],c_w_115);
AND_array_1506 AND_array_1506_i116(a,b[116],c_w_116);
AND_array_1506 AND_array_1506_i117(a,b[117],c_w_117);
AND_array_1506 AND_array_1506_i118(a,b[118],c_w_118);
AND_array_1506 AND_array_1506_i119(a,b[119],c_w_119);
AND_array_1506 AND_array_1506_i120(a,b[120],c_w_120);
AND_array_1506 AND_array_1506_i121(a,b[121],c_w_121);
AND_array_1506 AND_array_1506_i122(a,b[122],c_w_122);
AND_array_1506 AND_array_1506_i123(a,b[123],c_w_123);
AND_array_1506 AND_array_1506_i124(a,b[124],c_w_124);
AND_array_1506 AND_array_1506_i125(a,b[125],c_w_125);
AND_array_1506 AND_array_1506_i126(a,b[126],c_w_126);
AND_array_1506 AND_array_1506_i127(a,b[127],c_w_127);
AND_array_1506 AND_array_1506_i128(a,b[128],c_w_128);
AND_array_1506 AND_array_1506_i129(a,b[129],c_w_129);
AND_array_1506 AND_array_1506_i130(a,b[130],c_w_130);
AND_array_1506 AND_array_1506_i131(a,b[131],c_w_131);
AND_array_1506 AND_array_1506_i132(a,b[132],c_w_132);
AND_array_1506 AND_array_1506_i133(a,b[133],c_w_133);
AND_array_1506 AND_array_1506_i134(a,b[134],c_w_134);
AND_array_1506 AND_array_1506_i135(a,b[135],c_w_135);
AND_array_1506 AND_array_1506_i136(a,b[136],c_w_136);
AND_array_1506 AND_array_1506_i137(a,b[137],c_w_137);
AND_array_1506 AND_array_1506_i138(a,b[138],c_w_138);
AND_array_1506 AND_array_1506_i139(a,b[139],c_w_139);
AND_array_1506 AND_array_1506_i140(a,b[140],c_w_140);
AND_array_1506 AND_array_1506_i141(a,b[141],c_w_141);
AND_array_1506 AND_array_1506_i142(a,b[142],c_w_142);
AND_array_1506 AND_array_1506_i143(a,b[143],c_w_143);
AND_array_1506 AND_array_1506_i144(a,b[144],c_w_144);
AND_array_1506 AND_array_1506_i145(a,b[145],c_w_145);
AND_array_1506 AND_array_1506_i146(a,b[146],c_w_146);
AND_array_1506 AND_array_1506_i147(a,b[147],c_w_147);
AND_array_1506 AND_array_1506_i148(a,b[148],c_w_148);
AND_array_1506 AND_array_1506_i149(a,b[149],c_w_149);
AND_array_1506 AND_array_1506_i150(a,b[150],c_w_150);
AND_array_1506 AND_array_1506_i151(a,b[151],c_w_151);
AND_array_1506 AND_array_1506_i152(a,b[152],c_w_152);
AND_array_1506 AND_array_1506_i153(a,b[153],c_w_153);
AND_array_1506 AND_array_1506_i154(a,b[154],c_w_154);
AND_array_1506 AND_array_1506_i155(a,b[155],c_w_155);
AND_array_1506 AND_array_1506_i156(a,b[156],c_w_156);
AND_array_1506 AND_array_1506_i157(a,b[157],c_w_157);
AND_array_1506 AND_array_1506_i158(a,b[158],c_w_158);
AND_array_1506 AND_array_1506_i159(a,b[159],c_w_159);
AND_array_1506 AND_array_1506_i160(a,b[160],c_w_160);
AND_array_1506 AND_array_1506_i161(a,b[161],c_w_161);
AND_array_1506 AND_array_1506_i162(a,b[162],c_w_162);
AND_array_1506 AND_array_1506_i163(a,b[163],c_w_163);
AND_array_1506 AND_array_1506_i164(a,b[164],c_w_164);
AND_array_1506 AND_array_1506_i165(a,b[165],c_w_165);
AND_array_1506 AND_array_1506_i166(a,b[166],c_w_166);
AND_array_1506 AND_array_1506_i167(a,b[167],c_w_167);
AND_array_1506 AND_array_1506_i168(a,b[168],c_w_168);
AND_array_1506 AND_array_1506_i169(a,b[169],c_w_169);
AND_array_1506 AND_array_1506_i170(a,b[170],c_w_170);
AND_array_1506 AND_array_1506_i171(a,b[171],c_w_171);
AND_array_1506 AND_array_1506_i172(a,b[172],c_w_172);
AND_array_1506 AND_array_1506_i173(a,b[173],c_w_173);
AND_array_1506 AND_array_1506_i174(a,b[174],c_w_174);
AND_array_1506 AND_array_1506_i175(a,b[175],c_w_175);
AND_array_1506 AND_array_1506_i176(a,b[176],c_w_176);
AND_array_1506 AND_array_1506_i177(a,b[177],c_w_177);
AND_array_1506 AND_array_1506_i178(a,b[178],c_w_178);
AND_array_1506 AND_array_1506_i179(a,b[179],c_w_179);
AND_array_1506 AND_array_1506_i180(a,b[180],c_w_180);
AND_array_1506 AND_array_1506_i181(a,b[181],c_w_181);
AND_array_1506 AND_array_1506_i182(a,b[182],c_w_182);
AND_array_1506 AND_array_1506_i183(a,b[183],c_w_183);
AND_array_1506 AND_array_1506_i184(a,b[184],c_w_184);
AND_array_1506 AND_array_1506_i185(a,b[185],c_w_185);
AND_array_1506 AND_array_1506_i186(a,b[186],c_w_186);
AND_array_1506 AND_array_1506_i187(a,b[187],c_w_187);
AND_array_1506 AND_array_1506_i188(a,b[188],c_w_188);
AND_array_1506 AND_array_1506_i189(a,b[189],c_w_189);
AND_array_1506 AND_array_1506_i190(a,b[190],c_w_190);
AND_array_1506 AND_array_1506_i191(a,b[191],c_w_191);
AND_array_1506 AND_array_1506_i192(a,b[192],c_w_192);
AND_array_1506 AND_array_1506_i193(a,b[193],c_w_193);
AND_array_1506 AND_array_1506_i194(a,b[194],c_w_194);
AND_array_1506 AND_array_1506_i195(a,b[195],c_w_195);
AND_array_1506 AND_array_1506_i196(a,b[196],c_w_196);
AND_array_1506 AND_array_1506_i197(a,b[197],c_w_197);
AND_array_1506 AND_array_1506_i198(a,b[198],c_w_198);
AND_array_1506 AND_array_1506_i199(a,b[199],c_w_199);
AND_array_1506 AND_array_1506_i200(a,b[200],c_w_200);
AND_array_1506 AND_array_1506_i201(a,b[201],c_w_201);
AND_array_1506 AND_array_1506_i202(a,b[202],c_w_202);
AND_array_1506 AND_array_1506_i203(a,b[203],c_w_203);
AND_array_1506 AND_array_1506_i204(a,b[204],c_w_204);
AND_array_1506 AND_array_1506_i205(a,b[205],c_w_205);
AND_array_1506 AND_array_1506_i206(a,b[206],c_w_206);
AND_array_1506 AND_array_1506_i207(a,b[207],c_w_207);
AND_array_1506 AND_array_1506_i208(a,b[208],c_w_208);
AND_array_1506 AND_array_1506_i209(a,b[209],c_w_209);
AND_array_1506 AND_array_1506_i210(a,b[210],c_w_210);
AND_array_1506 AND_array_1506_i211(a,b[211],c_w_211);
AND_array_1506 AND_array_1506_i212(a,b[212],c_w_212);
AND_array_1506 AND_array_1506_i213(a,b[213],c_w_213);
AND_array_1506 AND_array_1506_i214(a,b[214],c_w_214);
AND_array_1506 AND_array_1506_i215(a,b[215],c_w_215);
AND_array_1506 AND_array_1506_i216(a,b[216],c_w_216);
AND_array_1506 AND_array_1506_i217(a,b[217],c_w_217);
AND_array_1506 AND_array_1506_i218(a,b[218],c_w_218);
AND_array_1506 AND_array_1506_i219(a,b[219],c_w_219);
AND_array_1506 AND_array_1506_i220(a,b[220],c_w_220);
AND_array_1506 AND_array_1506_i221(a,b[221],c_w_221);
AND_array_1506 AND_array_1506_i222(a,b[222],c_w_222);
AND_array_1506 AND_array_1506_i223(a,b[223],c_w_223);
AND_array_1506 AND_array_1506_i224(a,b[224],c_w_224);
AND_array_1506 AND_array_1506_i225(a,b[225],c_w_225);
AND_array_1506 AND_array_1506_i226(a,b[226],c_w_226);
AND_array_1506 AND_array_1506_i227(a,b[227],c_w_227);
AND_array_1506 AND_array_1506_i228(a,b[228],c_w_228);
AND_array_1506 AND_array_1506_i229(a,b[229],c_w_229);
AND_array_1506 AND_array_1506_i230(a,b[230],c_w_230);
AND_array_1506 AND_array_1506_i231(a,b[231],c_w_231);
AND_array_1506 AND_array_1506_i232(a,b[232],c_w_232);
AND_array_1506 AND_array_1506_i233(a,b[233],c_w_233);
AND_array_1506 AND_array_1506_i234(a,b[234],c_w_234);
AND_array_1506 AND_array_1506_i235(a,b[235],c_w_235);
AND_array_1506 AND_array_1506_i236(a,b[236],c_w_236);
AND_array_1506 AND_array_1506_i237(a,b[237],c_w_237);
AND_array_1506 AND_array_1506_i238(a,b[238],c_w_238);
AND_array_1506 AND_array_1506_i239(a,b[239],c_w_239);
AND_array_1506 AND_array_1506_i240(a,b[240],c_w_240);
AND_array_1506 AND_array_1506_i241(a,b[241],c_w_241);
AND_array_1506 AND_array_1506_i242(a,b[242],c_w_242);
AND_array_1506 AND_array_1506_i243(a,b[243],c_w_243);
AND_array_1506 AND_array_1506_i244(a,b[244],c_w_244);
AND_array_1506 AND_array_1506_i245(a,b[245],c_w_245);
AND_array_1506 AND_array_1506_i246(a,b[246],c_w_246);
AND_array_1506 AND_array_1506_i247(a,b[247],c_w_247);
AND_array_1506 AND_array_1506_i248(a,b[248],c_w_248);
AND_array_1506 AND_array_1506_i249(a,b[249],c_w_249);
AND_array_1506 AND_array_1506_i250(a,b[250],c_w_250);
AND_array_1506 AND_array_1506_i251(a,b[251],c_w_251);
AND_array_1506 AND_array_1506_i252(a,b[252],c_w_252);
AND_array_1506 AND_array_1506_i253(a,b[253],c_w_253);
AND_array_1506 AND_array_1506_i254(a,b[254],c_w_254);
AND_array_1506 AND_array_1506_i255(a,b[255],c_w_255);
AND_array_1506 AND_array_1506_i256(a,b[256],c_w_256);
AND_array_1506 AND_array_1506_i257(a,b[257],c_w_257);
AND_array_1506 AND_array_1506_i258(a,b[258],c_w_258);
AND_array_1506 AND_array_1506_i259(a,b[259],c_w_259);
AND_array_1506 AND_array_1506_i260(a,b[260],c_w_260);
AND_array_1506 AND_array_1506_i261(a,b[261],c_w_261);
AND_array_1506 AND_array_1506_i262(a,b[262],c_w_262);
AND_array_1506 AND_array_1506_i263(a,b[263],c_w_263);
AND_array_1506 AND_array_1506_i264(a,b[264],c_w_264);
AND_array_1506 AND_array_1506_i265(a,b[265],c_w_265);
AND_array_1506 AND_array_1506_i266(a,b[266],c_w_266);
AND_array_1506 AND_array_1506_i267(a,b[267],c_w_267);
AND_array_1506 AND_array_1506_i268(a,b[268],c_w_268);
AND_array_1506 AND_array_1506_i269(a,b[269],c_w_269);
AND_array_1506 AND_array_1506_i270(a,b[270],c_w_270);
AND_array_1506 AND_array_1506_i271(a,b[271],c_w_271);
AND_array_1506 AND_array_1506_i272(a,b[272],c_w_272);
AND_array_1506 AND_array_1506_i273(a,b[273],c_w_273);
AND_array_1506 AND_array_1506_i274(a,b[274],c_w_274);
AND_array_1506 AND_array_1506_i275(a,b[275],c_w_275);
AND_array_1506 AND_array_1506_i276(a,b[276],c_w_276);
AND_array_1506 AND_array_1506_i277(a,b[277],c_w_277);
AND_array_1506 AND_array_1506_i278(a,b[278],c_w_278);
AND_array_1506 AND_array_1506_i279(a,b[279],c_w_279);
AND_array_1506 AND_array_1506_i280(a,b[280],c_w_280);
AND_array_1506 AND_array_1506_i281(a,b[281],c_w_281);
AND_array_1506 AND_array_1506_i282(a,b[282],c_w_282);
AND_array_1506 AND_array_1506_i283(a,b[283],c_w_283);
AND_array_1506 AND_array_1506_i284(a,b[284],c_w_284);
AND_array_1506 AND_array_1506_i285(a,b[285],c_w_285);
AND_array_1506 AND_array_1506_i286(a,b[286],c_w_286);
AND_array_1506 AND_array_1506_i287(a,b[287],c_w_287);
AND_array_1506 AND_array_1506_i288(a,b[288],c_w_288);
AND_array_1506 AND_array_1506_i289(a,b[289],c_w_289);
AND_array_1506 AND_array_1506_i290(a,b[290],c_w_290);
AND_array_1506 AND_array_1506_i291(a,b[291],c_w_291);
AND_array_1506 AND_array_1506_i292(a,b[292],c_w_292);
AND_array_1506 AND_array_1506_i293(a,b[293],c_w_293);
AND_array_1506 AND_array_1506_i294(a,b[294],c_w_294);
AND_array_1506 AND_array_1506_i295(a,b[295],c_w_295);
AND_array_1506 AND_array_1506_i296(a,b[296],c_w_296);
AND_array_1506 AND_array_1506_i297(a,b[297],c_w_297);
AND_array_1506 AND_array_1506_i298(a,b[298],c_w_298);
AND_array_1506 AND_array_1506_i299(a,b[299],c_w_299);
AND_array_1506 AND_array_1506_i300(a,b[300],c_w_300);
AND_array_1506 AND_array_1506_i301(a,b[301],c_w_301);
AND_array_1506 AND_array_1506_i302(a,b[302],c_w_302);
AND_array_1506 AND_array_1506_i303(a,b[303],c_w_303);
AND_array_1506 AND_array_1506_i304(a,b[304],c_w_304);
AND_array_1506 AND_array_1506_i305(a,b[305],c_w_305);
AND_array_1506 AND_array_1506_i306(a,b[306],c_w_306);
AND_array_1506 AND_array_1506_i307(a,b[307],c_w_307);
AND_array_1506 AND_array_1506_i308(a,b[308],c_w_308);
AND_array_1506 AND_array_1506_i309(a,b[309],c_w_309);
AND_array_1506 AND_array_1506_i310(a,b[310],c_w_310);
AND_array_1506 AND_array_1506_i311(a,b[311],c_w_311);
AND_array_1506 AND_array_1506_i312(a,b[312],c_w_312);
AND_array_1506 AND_array_1506_i313(a,b[313],c_w_313);
AND_array_1506 AND_array_1506_i314(a,b[314],c_w_314);
AND_array_1506 AND_array_1506_i315(a,b[315],c_w_315);
AND_array_1506 AND_array_1506_i316(a,b[316],c_w_316);
AND_array_1506 AND_array_1506_i317(a,b[317],c_w_317);
AND_array_1506 AND_array_1506_i318(a,b[318],c_w_318);
AND_array_1506 AND_array_1506_i319(a,b[319],c_w_319);
AND_array_1506 AND_array_1506_i320(a,b[320],c_w_320);
AND_array_1506 AND_array_1506_i321(a,b[321],c_w_321);
AND_array_1506 AND_array_1506_i322(a,b[322],c_w_322);
AND_array_1506 AND_array_1506_i323(a,b[323],c_w_323);
AND_array_1506 AND_array_1506_i324(a,b[324],c_w_324);
AND_array_1506 AND_array_1506_i325(a,b[325],c_w_325);
AND_array_1506 AND_array_1506_i326(a,b[326],c_w_326);
AND_array_1506 AND_array_1506_i327(a,b[327],c_w_327);
AND_array_1506 AND_array_1506_i328(a,b[328],c_w_328);
AND_array_1506 AND_array_1506_i329(a,b[329],c_w_329);
AND_array_1506 AND_array_1506_i330(a,b[330],c_w_330);
AND_array_1506 AND_array_1506_i331(a,b[331],c_w_331);
AND_array_1506 AND_array_1506_i332(a,b[332],c_w_332);
AND_array_1506 AND_array_1506_i333(a,b[333],c_w_333);
AND_array_1506 AND_array_1506_i334(a,b[334],c_w_334);
AND_array_1506 AND_array_1506_i335(a,b[335],c_w_335);
AND_array_1506 AND_array_1506_i336(a,b[336],c_w_336);
AND_array_1506 AND_array_1506_i337(a,b[337],c_w_337);
AND_array_1506 AND_array_1506_i338(a,b[338],c_w_338);
AND_array_1506 AND_array_1506_i339(a,b[339],c_w_339);
AND_array_1506 AND_array_1506_i340(a,b[340],c_w_340);
AND_array_1506 AND_array_1506_i341(a,b[341],c_w_341);
AND_array_1506 AND_array_1506_i342(a,b[342],c_w_342);
AND_array_1506 AND_array_1506_i343(a,b[343],c_w_343);
AND_array_1506 AND_array_1506_i344(a,b[344],c_w_344);
AND_array_1506 AND_array_1506_i345(a,b[345],c_w_345);
AND_array_1506 AND_array_1506_i346(a,b[346],c_w_346);
AND_array_1506 AND_array_1506_i347(a,b[347],c_w_347);
AND_array_1506 AND_array_1506_i348(a,b[348],c_w_348);
AND_array_1506 AND_array_1506_i349(a,b[349],c_w_349);
AND_array_1506 AND_array_1506_i350(a,b[350],c_w_350);
AND_array_1506 AND_array_1506_i351(a,b[351],c_w_351);
AND_array_1506 AND_array_1506_i352(a,b[352],c_w_352);
AND_array_1506 AND_array_1506_i353(a,b[353],c_w_353);
AND_array_1506 AND_array_1506_i354(a,b[354],c_w_354);
AND_array_1506 AND_array_1506_i355(a,b[355],c_w_355);
AND_array_1506 AND_array_1506_i356(a,b[356],c_w_356);
AND_array_1506 AND_array_1506_i357(a,b[357],c_w_357);
AND_array_1506 AND_array_1506_i358(a,b[358],c_w_358);
AND_array_1506 AND_array_1506_i359(a,b[359],c_w_359);
AND_array_1506 AND_array_1506_i360(a,b[360],c_w_360);
AND_array_1506 AND_array_1506_i361(a,b[361],c_w_361);
AND_array_1506 AND_array_1506_i362(a,b[362],c_w_362);
AND_array_1506 AND_array_1506_i363(a,b[363],c_w_363);
AND_array_1506 AND_array_1506_i364(a,b[364],c_w_364);
AND_array_1506 AND_array_1506_i365(a,b[365],c_w_365);
AND_array_1506 AND_array_1506_i366(a,b[366],c_w_366);
AND_array_1506 AND_array_1506_i367(a,b[367],c_w_367);
AND_array_1506 AND_array_1506_i368(a,b[368],c_w_368);
AND_array_1506 AND_array_1506_i369(a,b[369],c_w_369);
AND_array_1506 AND_array_1506_i370(a,b[370],c_w_370);
AND_array_1506 AND_array_1506_i371(a,b[371],c_w_371);
AND_array_1506 AND_array_1506_i372(a,b[372],c_w_372);
AND_array_1506 AND_array_1506_i373(a,b[373],c_w_373);
AND_array_1506 AND_array_1506_i374(a,b[374],c_w_374);
AND_array_1506 AND_array_1506_i375(a,b[375],c_w_375);
AND_array_1506 AND_array_1506_i376(a,b[376],c_w_376);
AND_array_1506 AND_array_1506_i377(a,b[377],c_w_377);
AND_array_1506 AND_array_1506_i378(a,b[378],c_w_378);
AND_array_1506 AND_array_1506_i379(a,b[379],c_w_379);
AND_array_1506 AND_array_1506_i380(a,b[380],c_w_380);
AND_array_1506 AND_array_1506_i381(a,b[381],c_w_381);
AND_array_1506 AND_array_1506_i382(a,b[382],c_w_382);
AND_array_1506 AND_array_1506_i383(a,b[383],c_w_383);
AND_array_1506 AND_array_1506_i384(a,b[384],c_w_384);
AND_array_1506 AND_array_1506_i385(a,b[385],c_w_385);
AND_array_1506 AND_array_1506_i386(a,b[386],c_w_386);
AND_array_1506 AND_array_1506_i387(a,b[387],c_w_387);
AND_array_1506 AND_array_1506_i388(a,b[388],c_w_388);
AND_array_1506 AND_array_1506_i389(a,b[389],c_w_389);
AND_array_1506 AND_array_1506_i390(a,b[390],c_w_390);
AND_array_1506 AND_array_1506_i391(a,b[391],c_w_391);
AND_array_1506 AND_array_1506_i392(a,b[392],c_w_392);
AND_array_1506 AND_array_1506_i393(a,b[393],c_w_393);
AND_array_1506 AND_array_1506_i394(a,b[394],c_w_394);
AND_array_1506 AND_array_1506_i395(a,b[395],c_w_395);
AND_array_1506 AND_array_1506_i396(a,b[396],c_w_396);
AND_array_1506 AND_array_1506_i397(a,b[397],c_w_397);
AND_array_1506 AND_array_1506_i398(a,b[398],c_w_398);
AND_array_1506 AND_array_1506_i399(a,b[399],c_w_399);
AND_array_1506 AND_array_1506_i400(a,b[400],c_w_400);
AND_array_1506 AND_array_1506_i401(a,b[401],c_w_401);
AND_array_1506 AND_array_1506_i402(a,b[402],c_w_402);
AND_array_1506 AND_array_1506_i403(a,b[403],c_w_403);
AND_array_1506 AND_array_1506_i404(a,b[404],c_w_404);
AND_array_1506 AND_array_1506_i405(a,b[405],c_w_405);
AND_array_1506 AND_array_1506_i406(a,b[406],c_w_406);
AND_array_1506 AND_array_1506_i407(a,b[407],c_w_407);
AND_array_1506 AND_array_1506_i408(a,b[408],c_w_408);
AND_array_1506 AND_array_1506_i409(a,b[409],c_w_409);
AND_array_1506 AND_array_1506_i410(a,b[410],c_w_410);
AND_array_1506 AND_array_1506_i411(a,b[411],c_w_411);
AND_array_1506 AND_array_1506_i412(a,b[412],c_w_412);
AND_array_1506 AND_array_1506_i413(a,b[413],c_w_413);
AND_array_1506 AND_array_1506_i414(a,b[414],c_w_414);
AND_array_1506 AND_array_1506_i415(a,b[415],c_w_415);
AND_array_1506 AND_array_1506_i416(a,b[416],c_w_416);
AND_array_1506 AND_array_1506_i417(a,b[417],c_w_417);
AND_array_1506 AND_array_1506_i418(a,b[418],c_w_418);
AND_array_1506 AND_array_1506_i419(a,b[419],c_w_419);
AND_array_1506 AND_array_1506_i420(a,b[420],c_w_420);
AND_array_1506 AND_array_1506_i421(a,b[421],c_w_421);
AND_array_1506 AND_array_1506_i422(a,b[422],c_w_422);
AND_array_1506 AND_array_1506_i423(a,b[423],c_w_423);
AND_array_1506 AND_array_1506_i424(a,b[424],c_w_424);
AND_array_1506 AND_array_1506_i425(a,b[425],c_w_425);
AND_array_1506 AND_array_1506_i426(a,b[426],c_w_426);
AND_array_1506 AND_array_1506_i427(a,b[427],c_w_427);
AND_array_1506 AND_array_1506_i428(a,b[428],c_w_428);
AND_array_1506 AND_array_1506_i429(a,b[429],c_w_429);
AND_array_1506 AND_array_1506_i430(a,b[430],c_w_430);
AND_array_1506 AND_array_1506_i431(a,b[431],c_w_431);
AND_array_1506 AND_array_1506_i432(a,b[432],c_w_432);
AND_array_1506 AND_array_1506_i433(a,b[433],c_w_433);
AND_array_1506 AND_array_1506_i434(a,b[434],c_w_434);
AND_array_1506 AND_array_1506_i435(a,b[435],c_w_435);
AND_array_1506 AND_array_1506_i436(a,b[436],c_w_436);
AND_array_1506 AND_array_1506_i437(a,b[437],c_w_437);
AND_array_1506 AND_array_1506_i438(a,b[438],c_w_438);
AND_array_1506 AND_array_1506_i439(a,b[439],c_w_439);
AND_array_1506 AND_array_1506_i440(a,b[440],c_w_440);
AND_array_1506 AND_array_1506_i441(a,b[441],c_w_441);
AND_array_1506 AND_array_1506_i442(a,b[442],c_w_442);
AND_array_1506 AND_array_1506_i443(a,b[443],c_w_443);
AND_array_1506 AND_array_1506_i444(a,b[444],c_w_444);
AND_array_1506 AND_array_1506_i445(a,b[445],c_w_445);
AND_array_1506 AND_array_1506_i446(a,b[446],c_w_446);
AND_array_1506 AND_array_1506_i447(a,b[447],c_w_447);
AND_array_1506 AND_array_1506_i448(a,b[448],c_w_448);
AND_array_1506 AND_array_1506_i449(a,b[449],c_w_449);
AND_array_1506 AND_array_1506_i450(a,b[450],c_w_450);
AND_array_1506 AND_array_1506_i451(a,b[451],c_w_451);
AND_array_1506 AND_array_1506_i452(a,b[452],c_w_452);
AND_array_1506 AND_array_1506_i453(a,b[453],c_w_453);
AND_array_1506 AND_array_1506_i454(a,b[454],c_w_454);
AND_array_1506 AND_array_1506_i455(a,b[455],c_w_455);
AND_array_1506 AND_array_1506_i456(a,b[456],c_w_456);
AND_array_1506 AND_array_1506_i457(a,b[457],c_w_457);
AND_array_1506 AND_array_1506_i458(a,b[458],c_w_458);
AND_array_1506 AND_array_1506_i459(a,b[459],c_w_459);
AND_array_1506 AND_array_1506_i460(a,b[460],c_w_460);
AND_array_1506 AND_array_1506_i461(a,b[461],c_w_461);
AND_array_1506 AND_array_1506_i462(a,b[462],c_w_462);
AND_array_1506 AND_array_1506_i463(a,b[463],c_w_463);
AND_array_1506 AND_array_1506_i464(a,b[464],c_w_464);
AND_array_1506 AND_array_1506_i465(a,b[465],c_w_465);
AND_array_1506 AND_array_1506_i466(a,b[466],c_w_466);
AND_array_1506 AND_array_1506_i467(a,b[467],c_w_467);
AND_array_1506 AND_array_1506_i468(a,b[468],c_w_468);
AND_array_1506 AND_array_1506_i469(a,b[469],c_w_469);
AND_array_1506 AND_array_1506_i470(a,b[470],c_w_470);
AND_array_1506 AND_array_1506_i471(a,b[471],c_w_471);
AND_array_1506 AND_array_1506_i472(a,b[472],c_w_472);
AND_array_1506 AND_array_1506_i473(a,b[473],c_w_473);
AND_array_1506 AND_array_1506_i474(a,b[474],c_w_474);
AND_array_1506 AND_array_1506_i475(a,b[475],c_w_475);
AND_array_1506 AND_array_1506_i476(a,b[476],c_w_476);
AND_array_1506 AND_array_1506_i477(a,b[477],c_w_477);
AND_array_1506 AND_array_1506_i478(a,b[478],c_w_478);
AND_array_1506 AND_array_1506_i479(a,b[479],c_w_479);
AND_array_1506 AND_array_1506_i480(a,b[480],c_w_480);
AND_array_1506 AND_array_1506_i481(a,b[481],c_w_481);
AND_array_1506 AND_array_1506_i482(a,b[482],c_w_482);
AND_array_1506 AND_array_1506_i483(a,b[483],c_w_483);
AND_array_1506 AND_array_1506_i484(a,b[484],c_w_484);
AND_array_1506 AND_array_1506_i485(a,b[485],c_w_485);
AND_array_1506 AND_array_1506_i486(a,b[486],c_w_486);
AND_array_1506 AND_array_1506_i487(a,b[487],c_w_487);
AND_array_1506 AND_array_1506_i488(a,b[488],c_w_488);
AND_array_1506 AND_array_1506_i489(a,b[489],c_w_489);
AND_array_1506 AND_array_1506_i490(a,b[490],c_w_490);
AND_array_1506 AND_array_1506_i491(a,b[491],c_w_491);
AND_array_1506 AND_array_1506_i492(a,b[492],c_w_492);
AND_array_1506 AND_array_1506_i493(a,b[493],c_w_493);
AND_array_1506 AND_array_1506_i494(a,b[494],c_w_494);
AND_array_1506 AND_array_1506_i495(a,b[495],c_w_495);
AND_array_1506 AND_array_1506_i496(a,b[496],c_w_496);
AND_array_1506 AND_array_1506_i497(a,b[497],c_w_497);
AND_array_1506 AND_array_1506_i498(a,b[498],c_w_498);
AND_array_1506 AND_array_1506_i499(a,b[499],c_w_499);
AND_array_1506 AND_array_1506_i500(a,b[500],c_w_500);
AND_array_1506 AND_array_1506_i501(a,b[501],c_w_501);
AND_array_1506 AND_array_1506_i502(a,b[502],c_w_502);
AND_array_1506 AND_array_1506_i503(a,b[503],c_w_503);
AND_array_1506 AND_array_1506_i504(a,b[504],c_w_504);
AND_array_1506 AND_array_1506_i505(a,b[505],c_w_505);
AND_array_1506 AND_array_1506_i506(a,b[506],c_w_506);
AND_array_1506 AND_array_1506_i507(a,b[507],c_w_507);
AND_array_1506 AND_array_1506_i508(a,b[508],c_w_508);
AND_array_1506 AND_array_1506_i509(a,b[509],c_w_509);
AND_array_1506 AND_array_1506_i510(a,b[510],c_w_510);
AND_array_1506 AND_array_1506_i511(a,b[511],c_w_511);
AND_array_1506 AND_array_1506_i512(a,b[512],c_w_512);
AND_array_1506 AND_array_1506_i513(a,b[513],c_w_513);
AND_array_1506 AND_array_1506_i514(a,b[514],c_w_514);
AND_array_1506 AND_array_1506_i515(a,b[515],c_w_515);
AND_array_1506 AND_array_1506_i516(a,b[516],c_w_516);
AND_array_1506 AND_array_1506_i517(a,b[517],c_w_517);
AND_array_1506 AND_array_1506_i518(a,b[518],c_w_518);
AND_array_1506 AND_array_1506_i519(a,b[519],c_w_519);
AND_array_1506 AND_array_1506_i520(a,b[520],c_w_520);
AND_array_1506 AND_array_1506_i521(a,b[521],c_w_521);
AND_array_1506 AND_array_1506_i522(a,b[522],c_w_522);
AND_array_1506 AND_array_1506_i523(a,b[523],c_w_523);
AND_array_1506 AND_array_1506_i524(a,b[524],c_w_524);
AND_array_1506 AND_array_1506_i525(a,b[525],c_w_525);
AND_array_1506 AND_array_1506_i526(a,b[526],c_w_526);
AND_array_1506 AND_array_1506_i527(a,b[527],c_w_527);
AND_array_1506 AND_array_1506_i528(a,b[528],c_w_528);
AND_array_1506 AND_array_1506_i529(a,b[529],c_w_529);
AND_array_1506 AND_array_1506_i530(a,b[530],c_w_530);
AND_array_1506 AND_array_1506_i531(a,b[531],c_w_531);
AND_array_1506 AND_array_1506_i532(a,b[532],c_w_532);
AND_array_1506 AND_array_1506_i533(a,b[533],c_w_533);
AND_array_1506 AND_array_1506_i534(a,b[534],c_w_534);
AND_array_1506 AND_array_1506_i535(a,b[535],c_w_535);
AND_array_1506 AND_array_1506_i536(a,b[536],c_w_536);
AND_array_1506 AND_array_1506_i537(a,b[537],c_w_537);
AND_array_1506 AND_array_1506_i538(a,b[538],c_w_538);
AND_array_1506 AND_array_1506_i539(a,b[539],c_w_539);
AND_array_1506 AND_array_1506_i540(a,b[540],c_w_540);
AND_array_1506 AND_array_1506_i541(a,b[541],c_w_541);
AND_array_1506 AND_array_1506_i542(a,b[542],c_w_542);
AND_array_1506 AND_array_1506_i543(a,b[543],c_w_543);
AND_array_1506 AND_array_1506_i544(a,b[544],c_w_544);
AND_array_1506 AND_array_1506_i545(a,b[545],c_w_545);
AND_array_1506 AND_array_1506_i546(a,b[546],c_w_546);
AND_array_1506 AND_array_1506_i547(a,b[547],c_w_547);
AND_array_1506 AND_array_1506_i548(a,b[548],c_w_548);
AND_array_1506 AND_array_1506_i549(a,b[549],c_w_549);
AND_array_1506 AND_array_1506_i550(a,b[550],c_w_550);
AND_array_1506 AND_array_1506_i551(a,b[551],c_w_551);
AND_array_1506 AND_array_1506_i552(a,b[552],c_w_552);
AND_array_1506 AND_array_1506_i553(a,b[553],c_w_553);
AND_array_1506 AND_array_1506_i554(a,b[554],c_w_554);
AND_array_1506 AND_array_1506_i555(a,b[555],c_w_555);
AND_array_1506 AND_array_1506_i556(a,b[556],c_w_556);
AND_array_1506 AND_array_1506_i557(a,b[557],c_w_557);
AND_array_1506 AND_array_1506_i558(a,b[558],c_w_558);
AND_array_1506 AND_array_1506_i559(a,b[559],c_w_559);
AND_array_1506 AND_array_1506_i560(a,b[560],c_w_560);
AND_array_1506 AND_array_1506_i561(a,b[561],c_w_561);
AND_array_1506 AND_array_1506_i562(a,b[562],c_w_562);
AND_array_1506 AND_array_1506_i563(a,b[563],c_w_563);
AND_array_1506 AND_array_1506_i564(a,b[564],c_w_564);
AND_array_1506 AND_array_1506_i565(a,b[565],c_w_565);
AND_array_1506 AND_array_1506_i566(a,b[566],c_w_566);
AND_array_1506 AND_array_1506_i567(a,b[567],c_w_567);
AND_array_1506 AND_array_1506_i568(a,b[568],c_w_568);
AND_array_1506 AND_array_1506_i569(a,b[569],c_w_569);
AND_array_1506 AND_array_1506_i570(a,b[570],c_w_570);
AND_array_1506 AND_array_1506_i571(a,b[571],c_w_571);
AND_array_1506 AND_array_1506_i572(a,b[572],c_w_572);
AND_array_1506 AND_array_1506_i573(a,b[573],c_w_573);
AND_array_1506 AND_array_1506_i574(a,b[574],c_w_574);
AND_array_1506 AND_array_1506_i575(a,b[575],c_w_575);
AND_array_1506 AND_array_1506_i576(a,b[576],c_w_576);
AND_array_1506 AND_array_1506_i577(a,b[577],c_w_577);
AND_array_1506 AND_array_1506_i578(a,b[578],c_w_578);
AND_array_1506 AND_array_1506_i579(a,b[579],c_w_579);
AND_array_1506 AND_array_1506_i580(a,b[580],c_w_580);
AND_array_1506 AND_array_1506_i581(a,b[581],c_w_581);
AND_array_1506 AND_array_1506_i582(a,b[582],c_w_582);
AND_array_1506 AND_array_1506_i583(a,b[583],c_w_583);
AND_array_1506 AND_array_1506_i584(a,b[584],c_w_584);
AND_array_1506 AND_array_1506_i585(a,b[585],c_w_585);
AND_array_1506 AND_array_1506_i586(a,b[586],c_w_586);
AND_array_1506 AND_array_1506_i587(a,b[587],c_w_587);
AND_array_1506 AND_array_1506_i588(a,b[588],c_w_588);
AND_array_1506 AND_array_1506_i589(a,b[589],c_w_589);
AND_array_1506 AND_array_1506_i590(a,b[590],c_w_590);
AND_array_1506 AND_array_1506_i591(a,b[591],c_w_591);
AND_array_1506 AND_array_1506_i592(a,b[592],c_w_592);
AND_array_1506 AND_array_1506_i593(a,b[593],c_w_593);
AND_array_1506 AND_array_1506_i594(a,b[594],c_w_594);
AND_array_1506 AND_array_1506_i595(a,b[595],c_w_595);
AND_array_1506 AND_array_1506_i596(a,b[596],c_w_596);
AND_array_1506 AND_array_1506_i597(a,b[597],c_w_597);
AND_array_1506 AND_array_1506_i598(a,b[598],c_w_598);
AND_array_1506 AND_array_1506_i599(a,b[599],c_w_599);
AND_array_1506 AND_array_1506_i600(a,b[600],c_w_600);
AND_array_1506 AND_array_1506_i601(a,b[601],c_w_601);
AND_array_1506 AND_array_1506_i602(a,b[602],c_w_602);
AND_array_1506 AND_array_1506_i603(a,b[603],c_w_603);
AND_array_1506 AND_array_1506_i604(a,b[604],c_w_604);
AND_array_1506 AND_array_1506_i605(a,b[605],c_w_605);
AND_array_1506 AND_array_1506_i606(a,b[606],c_w_606);
AND_array_1506 AND_array_1506_i607(a,b[607],c_w_607);
AND_array_1506 AND_array_1506_i608(a,b[608],c_w_608);
AND_array_1506 AND_array_1506_i609(a,b[609],c_w_609);
AND_array_1506 AND_array_1506_i610(a,b[610],c_w_610);
AND_array_1506 AND_array_1506_i611(a,b[611],c_w_611);
AND_array_1506 AND_array_1506_i612(a,b[612],c_w_612);
AND_array_1506 AND_array_1506_i613(a,b[613],c_w_613);
AND_array_1506 AND_array_1506_i614(a,b[614],c_w_614);
AND_array_1506 AND_array_1506_i615(a,b[615],c_w_615);
AND_array_1506 AND_array_1506_i616(a,b[616],c_w_616);
AND_array_1506 AND_array_1506_i617(a,b[617],c_w_617);
AND_array_1506 AND_array_1506_i618(a,b[618],c_w_618);
AND_array_1506 AND_array_1506_i619(a,b[619],c_w_619);
AND_array_1506 AND_array_1506_i620(a,b[620],c_w_620);
AND_array_1506 AND_array_1506_i621(a,b[621],c_w_621);
AND_array_1506 AND_array_1506_i622(a,b[622],c_w_622);
AND_array_1506 AND_array_1506_i623(a,b[623],c_w_623);
AND_array_1506 AND_array_1506_i624(a,b[624],c_w_624);
AND_array_1506 AND_array_1506_i625(a,b[625],c_w_625);
AND_array_1506 AND_array_1506_i626(a,b[626],c_w_626);
AND_array_1506 AND_array_1506_i627(a,b[627],c_w_627);
AND_array_1506 AND_array_1506_i628(a,b[628],c_w_628);
AND_array_1506 AND_array_1506_i629(a,b[629],c_w_629);
AND_array_1506 AND_array_1506_i630(a,b[630],c_w_630);
AND_array_1506 AND_array_1506_i631(a,b[631],c_w_631);
AND_array_1506 AND_array_1506_i632(a,b[632],c_w_632);
AND_array_1506 AND_array_1506_i633(a,b[633],c_w_633);
AND_array_1506 AND_array_1506_i634(a,b[634],c_w_634);
AND_array_1506 AND_array_1506_i635(a,b[635],c_w_635);
AND_array_1506 AND_array_1506_i636(a,b[636],c_w_636);
AND_array_1506 AND_array_1506_i637(a,b[637],c_w_637);
AND_array_1506 AND_array_1506_i638(a,b[638],c_w_638);
AND_array_1506 AND_array_1506_i639(a,b[639],c_w_639);
AND_array_1506 AND_array_1506_i640(a,b[640],c_w_640);
AND_array_1506 AND_array_1506_i641(a,b[641],c_w_641);
AND_array_1506 AND_array_1506_i642(a,b[642],c_w_642);
AND_array_1506 AND_array_1506_i643(a,b[643],c_w_643);
AND_array_1506 AND_array_1506_i644(a,b[644],c_w_644);
AND_array_1506 AND_array_1506_i645(a,b[645],c_w_645);
AND_array_1506 AND_array_1506_i646(a,b[646],c_w_646);
AND_array_1506 AND_array_1506_i647(a,b[647],c_w_647);
AND_array_1506 AND_array_1506_i648(a,b[648],c_w_648);
AND_array_1506 AND_array_1506_i649(a,b[649],c_w_649);
AND_array_1506 AND_array_1506_i650(a,b[650],c_w_650);
AND_array_1506 AND_array_1506_i651(a,b[651],c_w_651);
AND_array_1506 AND_array_1506_i652(a,b[652],c_w_652);
AND_array_1506 AND_array_1506_i653(a,b[653],c_w_653);
AND_array_1506 AND_array_1506_i654(a,b[654],c_w_654);
AND_array_1506 AND_array_1506_i655(a,b[655],c_w_655);
AND_array_1506 AND_array_1506_i656(a,b[656],c_w_656);
AND_array_1506 AND_array_1506_i657(a,b[657],c_w_657);
AND_array_1506 AND_array_1506_i658(a,b[658],c_w_658);
AND_array_1506 AND_array_1506_i659(a,b[659],c_w_659);
AND_array_1506 AND_array_1506_i660(a,b[660],c_w_660);
AND_array_1506 AND_array_1506_i661(a,b[661],c_w_661);
AND_array_1506 AND_array_1506_i662(a,b[662],c_w_662);
AND_array_1506 AND_array_1506_i663(a,b[663],c_w_663);
AND_array_1506 AND_array_1506_i664(a,b[664],c_w_664);
AND_array_1506 AND_array_1506_i665(a,b[665],c_w_665);
AND_array_1506 AND_array_1506_i666(a,b[666],c_w_666);
AND_array_1506 AND_array_1506_i667(a,b[667],c_w_667);
AND_array_1506 AND_array_1506_i668(a,b[668],c_w_668);
AND_array_1506 AND_array_1506_i669(a,b[669],c_w_669);
AND_array_1506 AND_array_1506_i670(a,b[670],c_w_670);
AND_array_1506 AND_array_1506_i671(a,b[671],c_w_671);
AND_array_1506 AND_array_1506_i672(a,b[672],c_w_672);
AND_array_1506 AND_array_1506_i673(a,b[673],c_w_673);
AND_array_1506 AND_array_1506_i674(a,b[674],c_w_674);
AND_array_1506 AND_array_1506_i675(a,b[675],c_w_675);
AND_array_1506 AND_array_1506_i676(a,b[676],c_w_676);
AND_array_1506 AND_array_1506_i677(a,b[677],c_w_677);
AND_array_1506 AND_array_1506_i678(a,b[678],c_w_678);
AND_array_1506 AND_array_1506_i679(a,b[679],c_w_679);
AND_array_1506 AND_array_1506_i680(a,b[680],c_w_680);
AND_array_1506 AND_array_1506_i681(a,b[681],c_w_681);
AND_array_1506 AND_array_1506_i682(a,b[682],c_w_682);
AND_array_1506 AND_array_1506_i683(a,b[683],c_w_683);
AND_array_1506 AND_array_1506_i684(a,b[684],c_w_684);
AND_array_1506 AND_array_1506_i685(a,b[685],c_w_685);
AND_array_1506 AND_array_1506_i686(a,b[686],c_w_686);
AND_array_1506 AND_array_1506_i687(a,b[687],c_w_687);
AND_array_1506 AND_array_1506_i688(a,b[688],c_w_688);
AND_array_1506 AND_array_1506_i689(a,b[689],c_w_689);
AND_array_1506 AND_array_1506_i690(a,b[690],c_w_690);
AND_array_1506 AND_array_1506_i691(a,b[691],c_w_691);
AND_array_1506 AND_array_1506_i692(a,b[692],c_w_692);
AND_array_1506 AND_array_1506_i693(a,b[693],c_w_693);
AND_array_1506 AND_array_1506_i694(a,b[694],c_w_694);
AND_array_1506 AND_array_1506_i695(a,b[695],c_w_695);
AND_array_1506 AND_array_1506_i696(a,b[696],c_w_696);
AND_array_1506 AND_array_1506_i697(a,b[697],c_w_697);
AND_array_1506 AND_array_1506_i698(a,b[698],c_w_698);
AND_array_1506 AND_array_1506_i699(a,b[699],c_w_699);
AND_array_1506 AND_array_1506_i700(a,b[700],c_w_700);
AND_array_1506 AND_array_1506_i701(a,b[701],c_w_701);
AND_array_1506 AND_array_1506_i702(a,b[702],c_w_702);
AND_array_1506 AND_array_1506_i703(a,b[703],c_w_703);
AND_array_1506 AND_array_1506_i704(a,b[704],c_w_704);
AND_array_1506 AND_array_1506_i705(a,b[705],c_w_705);
AND_array_1506 AND_array_1506_i706(a,b[706],c_w_706);
AND_array_1506 AND_array_1506_i707(a,b[707],c_w_707);
AND_array_1506 AND_array_1506_i708(a,b[708],c_w_708);
AND_array_1506 AND_array_1506_i709(a,b[709],c_w_709);
AND_array_1506 AND_array_1506_i710(a,b[710],c_w_710);
AND_array_1506 AND_array_1506_i711(a,b[711],c_w_711);
AND_array_1506 AND_array_1506_i712(a,b[712],c_w_712);
AND_array_1506 AND_array_1506_i713(a,b[713],c_w_713);
AND_array_1506 AND_array_1506_i714(a,b[714],c_w_714);
AND_array_1506 AND_array_1506_i715(a,b[715],c_w_715);
AND_array_1506 AND_array_1506_i716(a,b[716],c_w_716);
AND_array_1506 AND_array_1506_i717(a,b[717],c_w_717);
AND_array_1506 AND_array_1506_i718(a,b[718],c_w_718);
AND_array_1506 AND_array_1506_i719(a,b[719],c_w_719);
AND_array_1506 AND_array_1506_i720(a,b[720],c_w_720);
AND_array_1506 AND_array_1506_i721(a,b[721],c_w_721);
AND_array_1506 AND_array_1506_i722(a,b[722],c_w_722);
AND_array_1506 AND_array_1506_i723(a,b[723],c_w_723);
AND_array_1506 AND_array_1506_i724(a,b[724],c_w_724);
AND_array_1506 AND_array_1506_i725(a,b[725],c_w_725);
AND_array_1506 AND_array_1506_i726(a,b[726],c_w_726);
AND_array_1506 AND_array_1506_i727(a,b[727],c_w_727);
AND_array_1506 AND_array_1506_i728(a,b[728],c_w_728);
AND_array_1506 AND_array_1506_i729(a,b[729],c_w_729);
AND_array_1506 AND_array_1506_i730(a,b[730],c_w_730);
AND_array_1506 AND_array_1506_i731(a,b[731],c_w_731);
AND_array_1506 AND_array_1506_i732(a,b[732],c_w_732);
AND_array_1506 AND_array_1506_i733(a,b[733],c_w_733);
AND_array_1506 AND_array_1506_i734(a,b[734],c_w_734);
AND_array_1506 AND_array_1506_i735(a,b[735],c_w_735);
AND_array_1506 AND_array_1506_i736(a,b[736],c_w_736);
AND_array_1506 AND_array_1506_i737(a,b[737],c_w_737);
AND_array_1506 AND_array_1506_i738(a,b[738],c_w_738);
AND_array_1506 AND_array_1506_i739(a,b[739],c_w_739);
AND_array_1506 AND_array_1506_i740(a,b[740],c_w_740);
AND_array_1506 AND_array_1506_i741(a,b[741],c_w_741);
AND_array_1506 AND_array_1506_i742(a,b[742],c_w_742);
AND_array_1506 AND_array_1506_i743(a,b[743],c_w_743);
AND_array_1506 AND_array_1506_i744(a,b[744],c_w_744);
AND_array_1506 AND_array_1506_i745(a,b[745],c_w_745);
AND_array_1506 AND_array_1506_i746(a,b[746],c_w_746);
AND_array_1506 AND_array_1506_i747(a,b[747],c_w_747);
AND_array_1506 AND_array_1506_i748(a,b[748],c_w_748);
AND_array_1506 AND_array_1506_i749(a,b[749],c_w_749);
AND_array_1506 AND_array_1506_i750(a,b[750],c_w_750);
AND_array_1506 AND_array_1506_i751(a,b[751],c_w_751);
AND_array_1506 AND_array_1506_i752(a,b[752],c_w_752);
AND_array_1506 AND_array_1506_i753(a,b[753],c_w_753);
AND_array_1506 AND_array_1506_i754(a,b[754],c_w_754);
AND_array_1506 AND_array_1506_i755(a,b[755],c_w_755);
AND_array_1506 AND_array_1506_i756(a,b[756],c_w_756);
AND_array_1506 AND_array_1506_i757(a,b[757],c_w_757);
AND_array_1506 AND_array_1506_i758(a,b[758],c_w_758);
AND_array_1506 AND_array_1506_i759(a,b[759],c_w_759);
AND_array_1506 AND_array_1506_i760(a,b[760],c_w_760);
AND_array_1506 AND_array_1506_i761(a,b[761],c_w_761);
AND_array_1506 AND_array_1506_i762(a,b[762],c_w_762);
AND_array_1506 AND_array_1506_i763(a,b[763],c_w_763);
AND_array_1506 AND_array_1506_i764(a,b[764],c_w_764);
AND_array_1506 AND_array_1506_i765(a,b[765],c_w_765);
AND_array_1506 AND_array_1506_i766(a,b[766],c_w_766);
AND_array_1506 AND_array_1506_i767(a,b[767],c_w_767);
AND_array_1506 AND_array_1506_i768(a,b[768],c_w_768);
AND_array_1506 AND_array_1506_i769(a,b[769],c_w_769);
AND_array_1506 AND_array_1506_i770(a,b[770],c_w_770);
AND_array_1506 AND_array_1506_i771(a,b[771],c_w_771);
AND_array_1506 AND_array_1506_i772(a,b[772],c_w_772);
AND_array_1506 AND_array_1506_i773(a,b[773],c_w_773);
AND_array_1506 AND_array_1506_i774(a,b[774],c_w_774);
AND_array_1506 AND_array_1506_i775(a,b[775],c_w_775);
AND_array_1506 AND_array_1506_i776(a,b[776],c_w_776);
AND_array_1506 AND_array_1506_i777(a,b[777],c_w_777);
AND_array_1506 AND_array_1506_i778(a,b[778],c_w_778);
AND_array_1506 AND_array_1506_i779(a,b[779],c_w_779);
AND_array_1506 AND_array_1506_i780(a,b[780],c_w_780);
AND_array_1506 AND_array_1506_i781(a,b[781],c_w_781);
AND_array_1506 AND_array_1506_i782(a,b[782],c_w_782);
AND_array_1506 AND_array_1506_i783(a,b[783],c_w_783);
AND_array_1506 AND_array_1506_i784(a,b[784],c_w_784);
AND_array_1506 AND_array_1506_i785(a,b[785],c_w_785);
AND_array_1506 AND_array_1506_i786(a,b[786],c_w_786);
AND_array_1506 AND_array_1506_i787(a,b[787],c_w_787);
AND_array_1506 AND_array_1506_i788(a,b[788],c_w_788);
AND_array_1506 AND_array_1506_i789(a,b[789],c_w_789);
AND_array_1506 AND_array_1506_i790(a,b[790],c_w_790);
AND_array_1506 AND_array_1506_i791(a,b[791],c_w_791);
AND_array_1506 AND_array_1506_i792(a,b[792],c_w_792);
AND_array_1506 AND_array_1506_i793(a,b[793],c_w_793);
AND_array_1506 AND_array_1506_i794(a,b[794],c_w_794);
AND_array_1506 AND_array_1506_i795(a,b[795],c_w_795);
AND_array_1506 AND_array_1506_i796(a,b[796],c_w_796);
AND_array_1506 AND_array_1506_i797(a,b[797],c_w_797);
AND_array_1506 AND_array_1506_i798(a,b[798],c_w_798);
AND_array_1506 AND_array_1506_i799(a,b[799],c_w_799);
AND_array_1506 AND_array_1506_i800(a,b[800],c_w_800);
AND_array_1506 AND_array_1506_i801(a,b[801],c_w_801);
AND_array_1506 AND_array_1506_i802(a,b[802],c_w_802);
AND_array_1506 AND_array_1506_i803(a,b[803],c_w_803);
AND_array_1506 AND_array_1506_i804(a,b[804],c_w_804);
AND_array_1506 AND_array_1506_i805(a,b[805],c_w_805);
AND_array_1506 AND_array_1506_i806(a,b[806],c_w_806);
AND_array_1506 AND_array_1506_i807(a,b[807],c_w_807);
AND_array_1506 AND_array_1506_i808(a,b[808],c_w_808);
AND_array_1506 AND_array_1506_i809(a,b[809],c_w_809);
AND_array_1506 AND_array_1506_i810(a,b[810],c_w_810);
AND_array_1506 AND_array_1506_i811(a,b[811],c_w_811);
AND_array_1506 AND_array_1506_i812(a,b[812],c_w_812);
AND_array_1506 AND_array_1506_i813(a,b[813],c_w_813);
AND_array_1506 AND_array_1506_i814(a,b[814],c_w_814);
AND_array_1506 AND_array_1506_i815(a,b[815],c_w_815);
AND_array_1506 AND_array_1506_i816(a,b[816],c_w_816);
AND_array_1506 AND_array_1506_i817(a,b[817],c_w_817);
AND_array_1506 AND_array_1506_i818(a,b[818],c_w_818);
AND_array_1506 AND_array_1506_i819(a,b[819],c_w_819);
AND_array_1506 AND_array_1506_i820(a,b[820],c_w_820);
AND_array_1506 AND_array_1506_i821(a,b[821],c_w_821);
AND_array_1506 AND_array_1506_i822(a,b[822],c_w_822);
AND_array_1506 AND_array_1506_i823(a,b[823],c_w_823);
AND_array_1506 AND_array_1506_i824(a,b[824],c_w_824);
AND_array_1506 AND_array_1506_i825(a,b[825],c_w_825);
AND_array_1506 AND_array_1506_i826(a,b[826],c_w_826);
AND_array_1506 AND_array_1506_i827(a,b[827],c_w_827);
AND_array_1506 AND_array_1506_i828(a,b[828],c_w_828);
AND_array_1506 AND_array_1506_i829(a,b[829],c_w_829);
AND_array_1506 AND_array_1506_i830(a,b[830],c_w_830);
AND_array_1506 AND_array_1506_i831(a,b[831],c_w_831);
AND_array_1506 AND_array_1506_i832(a,b[832],c_w_832);
AND_array_1506 AND_array_1506_i833(a,b[833],c_w_833);
AND_array_1506 AND_array_1506_i834(a,b[834],c_w_834);
AND_array_1506 AND_array_1506_i835(a,b[835],c_w_835);
AND_array_1506 AND_array_1506_i836(a,b[836],c_w_836);
AND_array_1506 AND_array_1506_i837(a,b[837],c_w_837);
AND_array_1506 AND_array_1506_i838(a,b[838],c_w_838);
AND_array_1506 AND_array_1506_i839(a,b[839],c_w_839);
AND_array_1506 AND_array_1506_i840(a,b[840],c_w_840);
AND_array_1506 AND_array_1506_i841(a,b[841],c_w_841);
AND_array_1506 AND_array_1506_i842(a,b[842],c_w_842);
AND_array_1506 AND_array_1506_i843(a,b[843],c_w_843);
AND_array_1506 AND_array_1506_i844(a,b[844],c_w_844);
AND_array_1506 AND_array_1506_i845(a,b[845],c_w_845);
AND_array_1506 AND_array_1506_i846(a,b[846],c_w_846);
AND_array_1506 AND_array_1506_i847(a,b[847],c_w_847);
AND_array_1506 AND_array_1506_i848(a,b[848],c_w_848);
AND_array_1506 AND_array_1506_i849(a,b[849],c_w_849);
AND_array_1506 AND_array_1506_i850(a,b[850],c_w_850);
AND_array_1506 AND_array_1506_i851(a,b[851],c_w_851);
AND_array_1506 AND_array_1506_i852(a,b[852],c_w_852);
AND_array_1506 AND_array_1506_i853(a,b[853],c_w_853);
AND_array_1506 AND_array_1506_i854(a,b[854],c_w_854);
AND_array_1506 AND_array_1506_i855(a,b[855],c_w_855);
AND_array_1506 AND_array_1506_i856(a,b[856],c_w_856);
AND_array_1506 AND_array_1506_i857(a,b[857],c_w_857);
AND_array_1506 AND_array_1506_i858(a,b[858],c_w_858);
AND_array_1506 AND_array_1506_i859(a,b[859],c_w_859);
AND_array_1506 AND_array_1506_i860(a,b[860],c_w_860);
AND_array_1506 AND_array_1506_i861(a,b[861],c_w_861);
AND_array_1506 AND_array_1506_i862(a,b[862],c_w_862);
AND_array_1506 AND_array_1506_i863(a,b[863],c_w_863);
AND_array_1506 AND_array_1506_i864(a,b[864],c_w_864);
AND_array_1506 AND_array_1506_i865(a,b[865],c_w_865);
AND_array_1506 AND_array_1506_i866(a,b[866],c_w_866);
AND_array_1506 AND_array_1506_i867(a,b[867],c_w_867);
AND_array_1506 AND_array_1506_i868(a,b[868],c_w_868);
AND_array_1506 AND_array_1506_i869(a,b[869],c_w_869);
AND_array_1506 AND_array_1506_i870(a,b[870],c_w_870);
AND_array_1506 AND_array_1506_i871(a,b[871],c_w_871);
AND_array_1506 AND_array_1506_i872(a,b[872],c_w_872);
AND_array_1506 AND_array_1506_i873(a,b[873],c_w_873);
AND_array_1506 AND_array_1506_i874(a,b[874],c_w_874);
AND_array_1506 AND_array_1506_i875(a,b[875],c_w_875);
AND_array_1506 AND_array_1506_i876(a,b[876],c_w_876);
AND_array_1506 AND_array_1506_i877(a,b[877],c_w_877);
AND_array_1506 AND_array_1506_i878(a,b[878],c_w_878);
AND_array_1506 AND_array_1506_i879(a,b[879],c_w_879);
AND_array_1506 AND_array_1506_i880(a,b[880],c_w_880);
AND_array_1506 AND_array_1506_i881(a,b[881],c_w_881);
AND_array_1506 AND_array_1506_i882(a,b[882],c_w_882);
AND_array_1506 AND_array_1506_i883(a,b[883],c_w_883);
AND_array_1506 AND_array_1506_i884(a,b[884],c_w_884);
AND_array_1506 AND_array_1506_i885(a,b[885],c_w_885);
AND_array_1506 AND_array_1506_i886(a,b[886],c_w_886);
AND_array_1506 AND_array_1506_i887(a,b[887],c_w_887);
AND_array_1506 AND_array_1506_i888(a,b[888],c_w_888);
AND_array_1506 AND_array_1506_i889(a,b[889],c_w_889);
AND_array_1506 AND_array_1506_i890(a,b[890],c_w_890);
AND_array_1506 AND_array_1506_i891(a,b[891],c_w_891);
AND_array_1506 AND_array_1506_i892(a,b[892],c_w_892);
AND_array_1506 AND_array_1506_i893(a,b[893],c_w_893);
AND_array_1506 AND_array_1506_i894(a,b[894],c_w_894);
AND_array_1506 AND_array_1506_i895(a,b[895],c_w_895);
AND_array_1506 AND_array_1506_i896(a,b[896],c_w_896);
AND_array_1506 AND_array_1506_i897(a,b[897],c_w_897);
AND_array_1506 AND_array_1506_i898(a,b[898],c_w_898);
AND_array_1506 AND_array_1506_i899(a,b[899],c_w_899);
AND_array_1506 AND_array_1506_i900(a,b[900],c_w_900);
AND_array_1506 AND_array_1506_i901(a,b[901],c_w_901);
AND_array_1506 AND_array_1506_i902(a,b[902],c_w_902);
AND_array_1506 AND_array_1506_i903(a,b[903],c_w_903);
AND_array_1506 AND_array_1506_i904(a,b[904],c_w_904);
AND_array_1506 AND_array_1506_i905(a,b[905],c_w_905);
AND_array_1506 AND_array_1506_i906(a,b[906],c_w_906);
AND_array_1506 AND_array_1506_i907(a,b[907],c_w_907);
AND_array_1506 AND_array_1506_i908(a,b[908],c_w_908);
AND_array_1506 AND_array_1506_i909(a,b[909],c_w_909);
AND_array_1506 AND_array_1506_i910(a,b[910],c_w_910);
AND_array_1506 AND_array_1506_i911(a,b[911],c_w_911);
AND_array_1506 AND_array_1506_i912(a,b[912],c_w_912);
AND_array_1506 AND_array_1506_i913(a,b[913],c_w_913);
AND_array_1506 AND_array_1506_i914(a,b[914],c_w_914);
AND_array_1506 AND_array_1506_i915(a,b[915],c_w_915);
AND_array_1506 AND_array_1506_i916(a,b[916],c_w_916);
AND_array_1506 AND_array_1506_i917(a,b[917],c_w_917);
AND_array_1506 AND_array_1506_i918(a,b[918],c_w_918);
AND_array_1506 AND_array_1506_i919(a,b[919],c_w_919);
AND_array_1506 AND_array_1506_i920(a,b[920],c_w_920);
AND_array_1506 AND_array_1506_i921(a,b[921],c_w_921);
AND_array_1506 AND_array_1506_i922(a,b[922],c_w_922);
AND_array_1506 AND_array_1506_i923(a,b[923],c_w_923);
AND_array_1506 AND_array_1506_i924(a,b[924],c_w_924);
AND_array_1506 AND_array_1506_i925(a,b[925],c_w_925);
AND_array_1506 AND_array_1506_i926(a,b[926],c_w_926);
AND_array_1506 AND_array_1506_i927(a,b[927],c_w_927);
AND_array_1506 AND_array_1506_i928(a,b[928],c_w_928);
AND_array_1506 AND_array_1506_i929(a,b[929],c_w_929);
AND_array_1506 AND_array_1506_i930(a,b[930],c_w_930);
AND_array_1506 AND_array_1506_i931(a,b[931],c_w_931);
AND_array_1506 AND_array_1506_i932(a,b[932],c_w_932);
AND_array_1506 AND_array_1506_i933(a,b[933],c_w_933);
AND_array_1506 AND_array_1506_i934(a,b[934],c_w_934);
AND_array_1506 AND_array_1506_i935(a,b[935],c_w_935);
AND_array_1506 AND_array_1506_i936(a,b[936],c_w_936);
AND_array_1506 AND_array_1506_i937(a,b[937],c_w_937);
AND_array_1506 AND_array_1506_i938(a,b[938],c_w_938);
AND_array_1506 AND_array_1506_i939(a,b[939],c_w_939);
AND_array_1506 AND_array_1506_i940(a,b[940],c_w_940);
AND_array_1506 AND_array_1506_i941(a,b[941],c_w_941);
AND_array_1506 AND_array_1506_i942(a,b[942],c_w_942);
AND_array_1506 AND_array_1506_i943(a,b[943],c_w_943);
AND_array_1506 AND_array_1506_i944(a,b[944],c_w_944);
AND_array_1506 AND_array_1506_i945(a,b[945],c_w_945);
AND_array_1506 AND_array_1506_i946(a,b[946],c_w_946);
AND_array_1506 AND_array_1506_i947(a,b[947],c_w_947);
AND_array_1506 AND_array_1506_i948(a,b[948],c_w_948);
AND_array_1506 AND_array_1506_i949(a,b[949],c_w_949);
AND_array_1506 AND_array_1506_i950(a,b[950],c_w_950);
AND_array_1506 AND_array_1506_i951(a,b[951],c_w_951);
AND_array_1506 AND_array_1506_i952(a,b[952],c_w_952);
AND_array_1506 AND_array_1506_i953(a,b[953],c_w_953);
AND_array_1506 AND_array_1506_i954(a,b[954],c_w_954);
AND_array_1506 AND_array_1506_i955(a,b[955],c_w_955);
AND_array_1506 AND_array_1506_i956(a,b[956],c_w_956);
AND_array_1506 AND_array_1506_i957(a,b[957],c_w_957);
AND_array_1506 AND_array_1506_i958(a,b[958],c_w_958);
AND_array_1506 AND_array_1506_i959(a,b[959],c_w_959);
AND_array_1506 AND_array_1506_i960(a,b[960],c_w_960);
AND_array_1506 AND_array_1506_i961(a,b[961],c_w_961);
AND_array_1506 AND_array_1506_i962(a,b[962],c_w_962);
AND_array_1506 AND_array_1506_i963(a,b[963],c_w_963);
AND_array_1506 AND_array_1506_i964(a,b[964],c_w_964);
AND_array_1506 AND_array_1506_i965(a,b[965],c_w_965);
AND_array_1506 AND_array_1506_i966(a,b[966],c_w_966);
AND_array_1506 AND_array_1506_i967(a,b[967],c_w_967);
AND_array_1506 AND_array_1506_i968(a,b[968],c_w_968);
AND_array_1506 AND_array_1506_i969(a,b[969],c_w_969);
AND_array_1506 AND_array_1506_i970(a,b[970],c_w_970);
AND_array_1506 AND_array_1506_i971(a,b[971],c_w_971);
AND_array_1506 AND_array_1506_i972(a,b[972],c_w_972);
AND_array_1506 AND_array_1506_i973(a,b[973],c_w_973);
AND_array_1506 AND_array_1506_i974(a,b[974],c_w_974);
AND_array_1506 AND_array_1506_i975(a,b[975],c_w_975);
AND_array_1506 AND_array_1506_i976(a,b[976],c_w_976);
AND_array_1506 AND_array_1506_i977(a,b[977],c_w_977);
AND_array_1506 AND_array_1506_i978(a,b[978],c_w_978);
AND_array_1506 AND_array_1506_i979(a,b[979],c_w_979);
AND_array_1506 AND_array_1506_i980(a,b[980],c_w_980);
AND_array_1506 AND_array_1506_i981(a,b[981],c_w_981);
AND_array_1506 AND_array_1506_i982(a,b[982],c_w_982);
AND_array_1506 AND_array_1506_i983(a,b[983],c_w_983);
AND_array_1506 AND_array_1506_i984(a,b[984],c_w_984);
AND_array_1506 AND_array_1506_i985(a,b[985],c_w_985);
AND_array_1506 AND_array_1506_i986(a,b[986],c_w_986);
AND_array_1506 AND_array_1506_i987(a,b[987],c_w_987);
AND_array_1506 AND_array_1506_i988(a,b[988],c_w_988);
AND_array_1506 AND_array_1506_i989(a,b[989],c_w_989);
AND_array_1506 AND_array_1506_i990(a,b[990],c_w_990);
AND_array_1506 AND_array_1506_i991(a,b[991],c_w_991);
AND_array_1506 AND_array_1506_i992(a,b[992],c_w_992);
AND_array_1506 AND_array_1506_i993(a,b[993],c_w_993);
AND_array_1506 AND_array_1506_i994(a,b[994],c_w_994);
AND_array_1506 AND_array_1506_i995(a,b[995],c_w_995);
AND_array_1506 AND_array_1506_i996(a,b[996],c_w_996);
AND_array_1506 AND_array_1506_i997(a,b[997],c_w_997);
AND_array_1506 AND_array_1506_i998(a,b[998],c_w_998);
AND_array_1506 AND_array_1506_i999(a,b[999],c_w_999);
AND_array_1506 AND_array_1506_i1000(a,b[1000],c_w_1000);
AND_array_1506 AND_array_1506_i1001(a,b[1001],c_w_1001);
AND_array_1506 AND_array_1506_i1002(a,b[1002],c_w_1002);
AND_array_1506 AND_array_1506_i1003(a,b[1003],c_w_1003);
AND_array_1506 AND_array_1506_i1004(a,b[1004],c_w_1004);
AND_array_1506 AND_array_1506_i1005(a,b[1005],c_w_1005);
AND_array_1506 AND_array_1506_i1006(a,b[1006],c_w_1006);
AND_array_1506 AND_array_1506_i1007(a,b[1007],c_w_1007);
AND_array_1506 AND_array_1506_i1008(a,b[1008],c_w_1008);
AND_array_1506 AND_array_1506_i1009(a,b[1009],c_w_1009);
AND_array_1506 AND_array_1506_i1010(a,b[1010],c_w_1010);
AND_array_1506 AND_array_1506_i1011(a,b[1011],c_w_1011);
AND_array_1506 AND_array_1506_i1012(a,b[1012],c_w_1012);
AND_array_1506 AND_array_1506_i1013(a,b[1013],c_w_1013);
AND_array_1506 AND_array_1506_i1014(a,b[1014],c_w_1014);
AND_array_1506 AND_array_1506_i1015(a,b[1015],c_w_1015);
AND_array_1506 AND_array_1506_i1016(a,b[1016],c_w_1016);
AND_array_1506 AND_array_1506_i1017(a,b[1017],c_w_1017);
AND_array_1506 AND_array_1506_i1018(a,b[1018],c_w_1018);
AND_array_1506 AND_array_1506_i1019(a,b[1019],c_w_1019);
AND_array_1506 AND_array_1506_i1020(a,b[1020],c_w_1020);
AND_array_1506 AND_array_1506_i1021(a,b[1021],c_w_1021);
AND_array_1506 AND_array_1506_i1022(a,b[1022],c_w_1022);
AND_array_1506 AND_array_1506_i1023(a,b[1023],c_w_1023);
AND_array_1506 AND_array_1506_i1024(a,b[1024],c_w_1024);
AND_array_1506 AND_array_1506_i1025(a,b[1025],c_w_1025);
AND_array_1506 AND_array_1506_i1026(a,b[1026],c_w_1026);
AND_array_1506 AND_array_1506_i1027(a,b[1027],c_w_1027);
AND_array_1506 AND_array_1506_i1028(a,b[1028],c_w_1028);
AND_array_1506 AND_array_1506_i1029(a,b[1029],c_w_1029);
AND_array_1506 AND_array_1506_i1030(a,b[1030],c_w_1030);
AND_array_1506 AND_array_1506_i1031(a,b[1031],c_w_1031);
AND_array_1506 AND_array_1506_i1032(a,b[1032],c_w_1032);
AND_array_1506 AND_array_1506_i1033(a,b[1033],c_w_1033);
AND_array_1506 AND_array_1506_i1034(a,b[1034],c_w_1034);
AND_array_1506 AND_array_1506_i1035(a,b[1035],c_w_1035);
AND_array_1506 AND_array_1506_i1036(a,b[1036],c_w_1036);
AND_array_1506 AND_array_1506_i1037(a,b[1037],c_w_1037);
AND_array_1506 AND_array_1506_i1038(a,b[1038],c_w_1038);
AND_array_1506 AND_array_1506_i1039(a,b[1039],c_w_1039);
AND_array_1506 AND_array_1506_i1040(a,b[1040],c_w_1040);
AND_array_1506 AND_array_1506_i1041(a,b[1041],c_w_1041);
AND_array_1506 AND_array_1506_i1042(a,b[1042],c_w_1042);
AND_array_1506 AND_array_1506_i1043(a,b[1043],c_w_1043);
AND_array_1506 AND_array_1506_i1044(a,b[1044],c_w_1044);
AND_array_1506 AND_array_1506_i1045(a,b[1045],c_w_1045);
AND_array_1506 AND_array_1506_i1046(a,b[1046],c_w_1046);
AND_array_1506 AND_array_1506_i1047(a,b[1047],c_w_1047);
AND_array_1506 AND_array_1506_i1048(a,b[1048],c_w_1048);
AND_array_1506 AND_array_1506_i1049(a,b[1049],c_w_1049);
AND_array_1506 AND_array_1506_i1050(a,b[1050],c_w_1050);
AND_array_1506 AND_array_1506_i1051(a,b[1051],c_w_1051);
AND_array_1506 AND_array_1506_i1052(a,b[1052],c_w_1052);
AND_array_1506 AND_array_1506_i1053(a,b[1053],c_w_1053);
AND_array_1506 AND_array_1506_i1054(a,b[1054],c_w_1054);
AND_array_1506 AND_array_1506_i1055(a,b[1055],c_w_1055);
AND_array_1506 AND_array_1506_i1056(a,b[1056],c_w_1056);
AND_array_1506 AND_array_1506_i1057(a,b[1057],c_w_1057);
AND_array_1506 AND_array_1506_i1058(a,b[1058],c_w_1058);
AND_array_1506 AND_array_1506_i1059(a,b[1059],c_w_1059);
AND_array_1506 AND_array_1506_i1060(a,b[1060],c_w_1060);
AND_array_1506 AND_array_1506_i1061(a,b[1061],c_w_1061);
AND_array_1506 AND_array_1506_i1062(a,b[1062],c_w_1062);
AND_array_1506 AND_array_1506_i1063(a,b[1063],c_w_1063);
AND_array_1506 AND_array_1506_i1064(a,b[1064],c_w_1064);
AND_array_1506 AND_array_1506_i1065(a,b[1065],c_w_1065);
AND_array_1506 AND_array_1506_i1066(a,b[1066],c_w_1066);
AND_array_1506 AND_array_1506_i1067(a,b[1067],c_w_1067);
AND_array_1506 AND_array_1506_i1068(a,b[1068],c_w_1068);
AND_array_1506 AND_array_1506_i1069(a,b[1069],c_w_1069);
AND_array_1506 AND_array_1506_i1070(a,b[1070],c_w_1070);
AND_array_1506 AND_array_1506_i1071(a,b[1071],c_w_1071);
AND_array_1506 AND_array_1506_i1072(a,b[1072],c_w_1072);
AND_array_1506 AND_array_1506_i1073(a,b[1073],c_w_1073);
AND_array_1506 AND_array_1506_i1074(a,b[1074],c_w_1074);
AND_array_1506 AND_array_1506_i1075(a,b[1075],c_w_1075);
AND_array_1506 AND_array_1506_i1076(a,b[1076],c_w_1076);
AND_array_1506 AND_array_1506_i1077(a,b[1077],c_w_1077);
AND_array_1506 AND_array_1506_i1078(a,b[1078],c_w_1078);
AND_array_1506 AND_array_1506_i1079(a,b[1079],c_w_1079);
AND_array_1506 AND_array_1506_i1080(a,b[1080],c_w_1080);
AND_array_1506 AND_array_1506_i1081(a,b[1081],c_w_1081);
AND_array_1506 AND_array_1506_i1082(a,b[1082],c_w_1082);
AND_array_1506 AND_array_1506_i1083(a,b[1083],c_w_1083);
AND_array_1506 AND_array_1506_i1084(a,b[1084],c_w_1084);
AND_array_1506 AND_array_1506_i1085(a,b[1085],c_w_1085);
AND_array_1506 AND_array_1506_i1086(a,b[1086],c_w_1086);
AND_array_1506 AND_array_1506_i1087(a,b[1087],c_w_1087);
AND_array_1506 AND_array_1506_i1088(a,b[1088],c_w_1088);
AND_array_1506 AND_array_1506_i1089(a,b[1089],c_w_1089);
AND_array_1506 AND_array_1506_i1090(a,b[1090],c_w_1090);
AND_array_1506 AND_array_1506_i1091(a,b[1091],c_w_1091);
AND_array_1506 AND_array_1506_i1092(a,b[1092],c_w_1092);
AND_array_1506 AND_array_1506_i1093(a,b[1093],c_w_1093);
AND_array_1506 AND_array_1506_i1094(a,b[1094],c_w_1094);
AND_array_1506 AND_array_1506_i1095(a,b[1095],c_w_1095);
AND_array_1506 AND_array_1506_i1096(a,b[1096],c_w_1096);
AND_array_1506 AND_array_1506_i1097(a,b[1097],c_w_1097);
AND_array_1506 AND_array_1506_i1098(a,b[1098],c_w_1098);
AND_array_1506 AND_array_1506_i1099(a,b[1099],c_w_1099);
AND_array_1506 AND_array_1506_i1100(a,b[1100],c_w_1100);
AND_array_1506 AND_array_1506_i1101(a,b[1101],c_w_1101);
AND_array_1506 AND_array_1506_i1102(a,b[1102],c_w_1102);
AND_array_1506 AND_array_1506_i1103(a,b[1103],c_w_1103);
AND_array_1506 AND_array_1506_i1104(a,b[1104],c_w_1104);
AND_array_1506 AND_array_1506_i1105(a,b[1105],c_w_1105);
AND_array_1506 AND_array_1506_i1106(a,b[1106],c_w_1106);
AND_array_1506 AND_array_1506_i1107(a,b[1107],c_w_1107);
AND_array_1506 AND_array_1506_i1108(a,b[1108],c_w_1108);
AND_array_1506 AND_array_1506_i1109(a,b[1109],c_w_1109);
AND_array_1506 AND_array_1506_i1110(a,b[1110],c_w_1110);
AND_array_1506 AND_array_1506_i1111(a,b[1111],c_w_1111);
AND_array_1506 AND_array_1506_i1112(a,b[1112],c_w_1112);
AND_array_1506 AND_array_1506_i1113(a,b[1113],c_w_1113);
AND_array_1506 AND_array_1506_i1114(a,b[1114],c_w_1114);
AND_array_1506 AND_array_1506_i1115(a,b[1115],c_w_1115);
AND_array_1506 AND_array_1506_i1116(a,b[1116],c_w_1116);
AND_array_1506 AND_array_1506_i1117(a,b[1117],c_w_1117);
AND_array_1506 AND_array_1506_i1118(a,b[1118],c_w_1118);
AND_array_1506 AND_array_1506_i1119(a,b[1119],c_w_1119);
AND_array_1506 AND_array_1506_i1120(a,b[1120],c_w_1120);
AND_array_1506 AND_array_1506_i1121(a,b[1121],c_w_1121);
AND_array_1506 AND_array_1506_i1122(a,b[1122],c_w_1122);
AND_array_1506 AND_array_1506_i1123(a,b[1123],c_w_1123);
AND_array_1506 AND_array_1506_i1124(a,b[1124],c_w_1124);
AND_array_1506 AND_array_1506_i1125(a,b[1125],c_w_1125);
AND_array_1506 AND_array_1506_i1126(a,b[1126],c_w_1126);
AND_array_1506 AND_array_1506_i1127(a,b[1127],c_w_1127);
AND_array_1506 AND_array_1506_i1128(a,b[1128],c_w_1128);
AND_array_1506 AND_array_1506_i1129(a,b[1129],c_w_1129);
AND_array_1506 AND_array_1506_i1130(a,b[1130],c_w_1130);
AND_array_1506 AND_array_1506_i1131(a,b[1131],c_w_1131);
AND_array_1506 AND_array_1506_i1132(a,b[1132],c_w_1132);
AND_array_1506 AND_array_1506_i1133(a,b[1133],c_w_1133);
AND_array_1506 AND_array_1506_i1134(a,b[1134],c_w_1134);
AND_array_1506 AND_array_1506_i1135(a,b[1135],c_w_1135);
AND_array_1506 AND_array_1506_i1136(a,b[1136],c_w_1136);
AND_array_1506 AND_array_1506_i1137(a,b[1137],c_w_1137);
AND_array_1506 AND_array_1506_i1138(a,b[1138],c_w_1138);
AND_array_1506 AND_array_1506_i1139(a,b[1139],c_w_1139);
AND_array_1506 AND_array_1506_i1140(a,b[1140],c_w_1140);
AND_array_1506 AND_array_1506_i1141(a,b[1141],c_w_1141);
AND_array_1506 AND_array_1506_i1142(a,b[1142],c_w_1142);
AND_array_1506 AND_array_1506_i1143(a,b[1143],c_w_1143);
AND_array_1506 AND_array_1506_i1144(a,b[1144],c_w_1144);
AND_array_1506 AND_array_1506_i1145(a,b[1145],c_w_1145);
AND_array_1506 AND_array_1506_i1146(a,b[1146],c_w_1146);
AND_array_1506 AND_array_1506_i1147(a,b[1147],c_w_1147);
AND_array_1506 AND_array_1506_i1148(a,b[1148],c_w_1148);
AND_array_1506 AND_array_1506_i1149(a,b[1149],c_w_1149);
AND_array_1506 AND_array_1506_i1150(a,b[1150],c_w_1150);
AND_array_1506 AND_array_1506_i1151(a,b[1151],c_w_1151);
AND_array_1506 AND_array_1506_i1152(a,b[1152],c_w_1152);
AND_array_1506 AND_array_1506_i1153(a,b[1153],c_w_1153);
AND_array_1506 AND_array_1506_i1154(a,b[1154],c_w_1154);
AND_array_1506 AND_array_1506_i1155(a,b[1155],c_w_1155);
AND_array_1506 AND_array_1506_i1156(a,b[1156],c_w_1156);
AND_array_1506 AND_array_1506_i1157(a,b[1157],c_w_1157);
AND_array_1506 AND_array_1506_i1158(a,b[1158],c_w_1158);
AND_array_1506 AND_array_1506_i1159(a,b[1159],c_w_1159);
AND_array_1506 AND_array_1506_i1160(a,b[1160],c_w_1160);
AND_array_1506 AND_array_1506_i1161(a,b[1161],c_w_1161);
AND_array_1506 AND_array_1506_i1162(a,b[1162],c_w_1162);
AND_array_1506 AND_array_1506_i1163(a,b[1163],c_w_1163);
AND_array_1506 AND_array_1506_i1164(a,b[1164],c_w_1164);
AND_array_1506 AND_array_1506_i1165(a,b[1165],c_w_1165);
AND_array_1506 AND_array_1506_i1166(a,b[1166],c_w_1166);
AND_array_1506 AND_array_1506_i1167(a,b[1167],c_w_1167);
AND_array_1506 AND_array_1506_i1168(a,b[1168],c_w_1168);
AND_array_1506 AND_array_1506_i1169(a,b[1169],c_w_1169);
AND_array_1506 AND_array_1506_i1170(a,b[1170],c_w_1170);
AND_array_1506 AND_array_1506_i1171(a,b[1171],c_w_1171);
AND_array_1506 AND_array_1506_i1172(a,b[1172],c_w_1172);
AND_array_1506 AND_array_1506_i1173(a,b[1173],c_w_1173);
AND_array_1506 AND_array_1506_i1174(a,b[1174],c_w_1174);
AND_array_1506 AND_array_1506_i1175(a,b[1175],c_w_1175);
AND_array_1506 AND_array_1506_i1176(a,b[1176],c_w_1176);
AND_array_1506 AND_array_1506_i1177(a,b[1177],c_w_1177);
AND_array_1506 AND_array_1506_i1178(a,b[1178],c_w_1178);
AND_array_1506 AND_array_1506_i1179(a,b[1179],c_w_1179);
AND_array_1506 AND_array_1506_i1180(a,b[1180],c_w_1180);
AND_array_1506 AND_array_1506_i1181(a,b[1181],c_w_1181);
AND_array_1506 AND_array_1506_i1182(a,b[1182],c_w_1182);
AND_array_1506 AND_array_1506_i1183(a,b[1183],c_w_1183);
AND_array_1506 AND_array_1506_i1184(a,b[1184],c_w_1184);
AND_array_1506 AND_array_1506_i1185(a,b[1185],c_w_1185);
AND_array_1506 AND_array_1506_i1186(a,b[1186],c_w_1186);
AND_array_1506 AND_array_1506_i1187(a,b[1187],c_w_1187);
AND_array_1506 AND_array_1506_i1188(a,b[1188],c_w_1188);
AND_array_1506 AND_array_1506_i1189(a,b[1189],c_w_1189);
AND_array_1506 AND_array_1506_i1190(a,b[1190],c_w_1190);
AND_array_1506 AND_array_1506_i1191(a,b[1191],c_w_1191);
AND_array_1506 AND_array_1506_i1192(a,b[1192],c_w_1192);
AND_array_1506 AND_array_1506_i1193(a,b[1193],c_w_1193);
AND_array_1506 AND_array_1506_i1194(a,b[1194],c_w_1194);
AND_array_1506 AND_array_1506_i1195(a,b[1195],c_w_1195);
AND_array_1506 AND_array_1506_i1196(a,b[1196],c_w_1196);
AND_array_1506 AND_array_1506_i1197(a,b[1197],c_w_1197);
AND_array_1506 AND_array_1506_i1198(a,b[1198],c_w_1198);
AND_array_1506 AND_array_1506_i1199(a,b[1199],c_w_1199);
AND_array_1506 AND_array_1506_i1200(a,b[1200],c_w_1200);
AND_array_1506 AND_array_1506_i1201(a,b[1201],c_w_1201);
AND_array_1506 AND_array_1506_i1202(a,b[1202],c_w_1202);
AND_array_1506 AND_array_1506_i1203(a,b[1203],c_w_1203);
AND_array_1506 AND_array_1506_i1204(a,b[1204],c_w_1204);
AND_array_1506 AND_array_1506_i1205(a,b[1205],c_w_1205);
AND_array_1506 AND_array_1506_i1206(a,b[1206],c_w_1206);
AND_array_1506 AND_array_1506_i1207(a,b[1207],c_w_1207);
AND_array_1506 AND_array_1506_i1208(a,b[1208],c_w_1208);
AND_array_1506 AND_array_1506_i1209(a,b[1209],c_w_1209);
AND_array_1506 AND_array_1506_i1210(a,b[1210],c_w_1210);
AND_array_1506 AND_array_1506_i1211(a,b[1211],c_w_1211);
AND_array_1506 AND_array_1506_i1212(a,b[1212],c_w_1212);
AND_array_1506 AND_array_1506_i1213(a,b[1213],c_w_1213);
AND_array_1506 AND_array_1506_i1214(a,b[1214],c_w_1214);
AND_array_1506 AND_array_1506_i1215(a,b[1215],c_w_1215);
AND_array_1506 AND_array_1506_i1216(a,b[1216],c_w_1216);
AND_array_1506 AND_array_1506_i1217(a,b[1217],c_w_1217);
AND_array_1506 AND_array_1506_i1218(a,b[1218],c_w_1218);
AND_array_1506 AND_array_1506_i1219(a,b[1219],c_w_1219);
AND_array_1506 AND_array_1506_i1220(a,b[1220],c_w_1220);
AND_array_1506 AND_array_1506_i1221(a,b[1221],c_w_1221);
AND_array_1506 AND_array_1506_i1222(a,b[1222],c_w_1222);
AND_array_1506 AND_array_1506_i1223(a,b[1223],c_w_1223);
AND_array_1506 AND_array_1506_i1224(a,b[1224],c_w_1224);
AND_array_1506 AND_array_1506_i1225(a,b[1225],c_w_1225);
AND_array_1506 AND_array_1506_i1226(a,b[1226],c_w_1226);
AND_array_1506 AND_array_1506_i1227(a,b[1227],c_w_1227);
AND_array_1506 AND_array_1506_i1228(a,b[1228],c_w_1228);
AND_array_1506 AND_array_1506_i1229(a,b[1229],c_w_1229);
AND_array_1506 AND_array_1506_i1230(a,b[1230],c_w_1230);
AND_array_1506 AND_array_1506_i1231(a,b[1231],c_w_1231);
AND_array_1506 AND_array_1506_i1232(a,b[1232],c_w_1232);
AND_array_1506 AND_array_1506_i1233(a,b[1233],c_w_1233);
AND_array_1506 AND_array_1506_i1234(a,b[1234],c_w_1234);
AND_array_1506 AND_array_1506_i1235(a,b[1235],c_w_1235);
AND_array_1506 AND_array_1506_i1236(a,b[1236],c_w_1236);
AND_array_1506 AND_array_1506_i1237(a,b[1237],c_w_1237);
AND_array_1506 AND_array_1506_i1238(a,b[1238],c_w_1238);
AND_array_1506 AND_array_1506_i1239(a,b[1239],c_w_1239);
AND_array_1506 AND_array_1506_i1240(a,b[1240],c_w_1240);
AND_array_1506 AND_array_1506_i1241(a,b[1241],c_w_1241);
AND_array_1506 AND_array_1506_i1242(a,b[1242],c_w_1242);
AND_array_1506 AND_array_1506_i1243(a,b[1243],c_w_1243);
AND_array_1506 AND_array_1506_i1244(a,b[1244],c_w_1244);
AND_array_1506 AND_array_1506_i1245(a,b[1245],c_w_1245);
AND_array_1506 AND_array_1506_i1246(a,b[1246],c_w_1246);
AND_array_1506 AND_array_1506_i1247(a,b[1247],c_w_1247);
AND_array_1506 AND_array_1506_i1248(a,b[1248],c_w_1248);
AND_array_1506 AND_array_1506_i1249(a,b[1249],c_w_1249);
AND_array_1506 AND_array_1506_i1250(a,b[1250],c_w_1250);
AND_array_1506 AND_array_1506_i1251(a,b[1251],c_w_1251);
AND_array_1506 AND_array_1506_i1252(a,b[1252],c_w_1252);
AND_array_1506 AND_array_1506_i1253(a,b[1253],c_w_1253);
AND_array_1506 AND_array_1506_i1254(a,b[1254],c_w_1254);
AND_array_1506 AND_array_1506_i1255(a,b[1255],c_w_1255);
AND_array_1506 AND_array_1506_i1256(a,b[1256],c_w_1256);
AND_array_1506 AND_array_1506_i1257(a,b[1257],c_w_1257);
AND_array_1506 AND_array_1506_i1258(a,b[1258],c_w_1258);
AND_array_1506 AND_array_1506_i1259(a,b[1259],c_w_1259);
AND_array_1506 AND_array_1506_i1260(a,b[1260],c_w_1260);
AND_array_1506 AND_array_1506_i1261(a,b[1261],c_w_1261);
AND_array_1506 AND_array_1506_i1262(a,b[1262],c_w_1262);
AND_array_1506 AND_array_1506_i1263(a,b[1263],c_w_1263);
AND_array_1506 AND_array_1506_i1264(a,b[1264],c_w_1264);
AND_array_1506 AND_array_1506_i1265(a,b[1265],c_w_1265);
AND_array_1506 AND_array_1506_i1266(a,b[1266],c_w_1266);
AND_array_1506 AND_array_1506_i1267(a,b[1267],c_w_1267);
AND_array_1506 AND_array_1506_i1268(a,b[1268],c_w_1268);
AND_array_1506 AND_array_1506_i1269(a,b[1269],c_w_1269);
AND_array_1506 AND_array_1506_i1270(a,b[1270],c_w_1270);
AND_array_1506 AND_array_1506_i1271(a,b[1271],c_w_1271);
AND_array_1506 AND_array_1506_i1272(a,b[1272],c_w_1272);
AND_array_1506 AND_array_1506_i1273(a,b[1273],c_w_1273);
AND_array_1506 AND_array_1506_i1274(a,b[1274],c_w_1274);
AND_array_1506 AND_array_1506_i1275(a,b[1275],c_w_1275);
AND_array_1506 AND_array_1506_i1276(a,b[1276],c_w_1276);
AND_array_1506 AND_array_1506_i1277(a,b[1277],c_w_1277);
AND_array_1506 AND_array_1506_i1278(a,b[1278],c_w_1278);
AND_array_1506 AND_array_1506_i1279(a,b[1279],c_w_1279);
AND_array_1506 AND_array_1506_i1280(a,b[1280],c_w_1280);
AND_array_1506 AND_array_1506_i1281(a,b[1281],c_w_1281);
AND_array_1506 AND_array_1506_i1282(a,b[1282],c_w_1282);
AND_array_1506 AND_array_1506_i1283(a,b[1283],c_w_1283);
AND_array_1506 AND_array_1506_i1284(a,b[1284],c_w_1284);
AND_array_1506 AND_array_1506_i1285(a,b[1285],c_w_1285);
AND_array_1506 AND_array_1506_i1286(a,b[1286],c_w_1286);
AND_array_1506 AND_array_1506_i1287(a,b[1287],c_w_1287);
AND_array_1506 AND_array_1506_i1288(a,b[1288],c_w_1288);
AND_array_1506 AND_array_1506_i1289(a,b[1289],c_w_1289);
AND_array_1506 AND_array_1506_i1290(a,b[1290],c_w_1290);
AND_array_1506 AND_array_1506_i1291(a,b[1291],c_w_1291);
AND_array_1506 AND_array_1506_i1292(a,b[1292],c_w_1292);
AND_array_1506 AND_array_1506_i1293(a,b[1293],c_w_1293);
AND_array_1506 AND_array_1506_i1294(a,b[1294],c_w_1294);
AND_array_1506 AND_array_1506_i1295(a,b[1295],c_w_1295);
AND_array_1506 AND_array_1506_i1296(a,b[1296],c_w_1296);
AND_array_1506 AND_array_1506_i1297(a,b[1297],c_w_1297);
AND_array_1506 AND_array_1506_i1298(a,b[1298],c_w_1298);
AND_array_1506 AND_array_1506_i1299(a,b[1299],c_w_1299);
AND_array_1506 AND_array_1506_i1300(a,b[1300],c_w_1300);
AND_array_1506 AND_array_1506_i1301(a,b[1301],c_w_1301);
AND_array_1506 AND_array_1506_i1302(a,b[1302],c_w_1302);
AND_array_1506 AND_array_1506_i1303(a,b[1303],c_w_1303);
AND_array_1506 AND_array_1506_i1304(a,b[1304],c_w_1304);
AND_array_1506 AND_array_1506_i1305(a,b[1305],c_w_1305);
AND_array_1506 AND_array_1506_i1306(a,b[1306],c_w_1306);
AND_array_1506 AND_array_1506_i1307(a,b[1307],c_w_1307);
AND_array_1506 AND_array_1506_i1308(a,b[1308],c_w_1308);
AND_array_1506 AND_array_1506_i1309(a,b[1309],c_w_1309);
AND_array_1506 AND_array_1506_i1310(a,b[1310],c_w_1310);
AND_array_1506 AND_array_1506_i1311(a,b[1311],c_w_1311);
AND_array_1506 AND_array_1506_i1312(a,b[1312],c_w_1312);
AND_array_1506 AND_array_1506_i1313(a,b[1313],c_w_1313);
AND_array_1506 AND_array_1506_i1314(a,b[1314],c_w_1314);
AND_array_1506 AND_array_1506_i1315(a,b[1315],c_w_1315);
AND_array_1506 AND_array_1506_i1316(a,b[1316],c_w_1316);
AND_array_1506 AND_array_1506_i1317(a,b[1317],c_w_1317);
AND_array_1506 AND_array_1506_i1318(a,b[1318],c_w_1318);
AND_array_1506 AND_array_1506_i1319(a,b[1319],c_w_1319);
AND_array_1506 AND_array_1506_i1320(a,b[1320],c_w_1320);
AND_array_1506 AND_array_1506_i1321(a,b[1321],c_w_1321);
AND_array_1506 AND_array_1506_i1322(a,b[1322],c_w_1322);
AND_array_1506 AND_array_1506_i1323(a,b[1323],c_w_1323);
AND_array_1506 AND_array_1506_i1324(a,b[1324],c_w_1324);
AND_array_1506 AND_array_1506_i1325(a,b[1325],c_w_1325);
AND_array_1506 AND_array_1506_i1326(a,b[1326],c_w_1326);
AND_array_1506 AND_array_1506_i1327(a,b[1327],c_w_1327);
AND_array_1506 AND_array_1506_i1328(a,b[1328],c_w_1328);
AND_array_1506 AND_array_1506_i1329(a,b[1329],c_w_1329);
AND_array_1506 AND_array_1506_i1330(a,b[1330],c_w_1330);
AND_array_1506 AND_array_1506_i1331(a,b[1331],c_w_1331);
AND_array_1506 AND_array_1506_i1332(a,b[1332],c_w_1332);
AND_array_1506 AND_array_1506_i1333(a,b[1333],c_w_1333);
AND_array_1506 AND_array_1506_i1334(a,b[1334],c_w_1334);
AND_array_1506 AND_array_1506_i1335(a,b[1335],c_w_1335);
AND_array_1506 AND_array_1506_i1336(a,b[1336],c_w_1336);
AND_array_1506 AND_array_1506_i1337(a,b[1337],c_w_1337);
AND_array_1506 AND_array_1506_i1338(a,b[1338],c_w_1338);
AND_array_1506 AND_array_1506_i1339(a,b[1339],c_w_1339);
AND_array_1506 AND_array_1506_i1340(a,b[1340],c_w_1340);
AND_array_1506 AND_array_1506_i1341(a,b[1341],c_w_1341);
AND_array_1506 AND_array_1506_i1342(a,b[1342],c_w_1342);
AND_array_1506 AND_array_1506_i1343(a,b[1343],c_w_1343);
AND_array_1506 AND_array_1506_i1344(a,b[1344],c_w_1344);
AND_array_1506 AND_array_1506_i1345(a,b[1345],c_w_1345);
AND_array_1506 AND_array_1506_i1346(a,b[1346],c_w_1346);
AND_array_1506 AND_array_1506_i1347(a,b[1347],c_w_1347);
AND_array_1506 AND_array_1506_i1348(a,b[1348],c_w_1348);
AND_array_1506 AND_array_1506_i1349(a,b[1349],c_w_1349);
AND_array_1506 AND_array_1506_i1350(a,b[1350],c_w_1350);
AND_array_1506 AND_array_1506_i1351(a,b[1351],c_w_1351);
AND_array_1506 AND_array_1506_i1352(a,b[1352],c_w_1352);
AND_array_1506 AND_array_1506_i1353(a,b[1353],c_w_1353);
AND_array_1506 AND_array_1506_i1354(a,b[1354],c_w_1354);
AND_array_1506 AND_array_1506_i1355(a,b[1355],c_w_1355);
AND_array_1506 AND_array_1506_i1356(a,b[1356],c_w_1356);
AND_array_1506 AND_array_1506_i1357(a,b[1357],c_w_1357);
AND_array_1506 AND_array_1506_i1358(a,b[1358],c_w_1358);
AND_array_1506 AND_array_1506_i1359(a,b[1359],c_w_1359);
AND_array_1506 AND_array_1506_i1360(a,b[1360],c_w_1360);
AND_array_1506 AND_array_1506_i1361(a,b[1361],c_w_1361);
AND_array_1506 AND_array_1506_i1362(a,b[1362],c_w_1362);
AND_array_1506 AND_array_1506_i1363(a,b[1363],c_w_1363);
AND_array_1506 AND_array_1506_i1364(a,b[1364],c_w_1364);
AND_array_1506 AND_array_1506_i1365(a,b[1365],c_w_1365);
AND_array_1506 AND_array_1506_i1366(a,b[1366],c_w_1366);
AND_array_1506 AND_array_1506_i1367(a,b[1367],c_w_1367);
AND_array_1506 AND_array_1506_i1368(a,b[1368],c_w_1368);
AND_array_1506 AND_array_1506_i1369(a,b[1369],c_w_1369);
AND_array_1506 AND_array_1506_i1370(a,b[1370],c_w_1370);
AND_array_1506 AND_array_1506_i1371(a,b[1371],c_w_1371);
AND_array_1506 AND_array_1506_i1372(a,b[1372],c_w_1372);
AND_array_1506 AND_array_1506_i1373(a,b[1373],c_w_1373);
AND_array_1506 AND_array_1506_i1374(a,b[1374],c_w_1374);
AND_array_1506 AND_array_1506_i1375(a,b[1375],c_w_1375);
AND_array_1506 AND_array_1506_i1376(a,b[1376],c_w_1376);
AND_array_1506 AND_array_1506_i1377(a,b[1377],c_w_1377);
AND_array_1506 AND_array_1506_i1378(a,b[1378],c_w_1378);
AND_array_1506 AND_array_1506_i1379(a,b[1379],c_w_1379);
AND_array_1506 AND_array_1506_i1380(a,b[1380],c_w_1380);
AND_array_1506 AND_array_1506_i1381(a,b[1381],c_w_1381);
AND_array_1506 AND_array_1506_i1382(a,b[1382],c_w_1382);
AND_array_1506 AND_array_1506_i1383(a,b[1383],c_w_1383);
AND_array_1506 AND_array_1506_i1384(a,b[1384],c_w_1384);
AND_array_1506 AND_array_1506_i1385(a,b[1385],c_w_1385);
AND_array_1506 AND_array_1506_i1386(a,b[1386],c_w_1386);
AND_array_1506 AND_array_1506_i1387(a,b[1387],c_w_1387);
AND_array_1506 AND_array_1506_i1388(a,b[1388],c_w_1388);
AND_array_1506 AND_array_1506_i1389(a,b[1389],c_w_1389);
AND_array_1506 AND_array_1506_i1390(a,b[1390],c_w_1390);
AND_array_1506 AND_array_1506_i1391(a,b[1391],c_w_1391);
AND_array_1506 AND_array_1506_i1392(a,b[1392],c_w_1392);
AND_array_1506 AND_array_1506_i1393(a,b[1393],c_w_1393);
AND_array_1506 AND_array_1506_i1394(a,b[1394],c_w_1394);
AND_array_1506 AND_array_1506_i1395(a,b[1395],c_w_1395);
AND_array_1506 AND_array_1506_i1396(a,b[1396],c_w_1396);
AND_array_1506 AND_array_1506_i1397(a,b[1397],c_w_1397);
AND_array_1506 AND_array_1506_i1398(a,b[1398],c_w_1398);
AND_array_1506 AND_array_1506_i1399(a,b[1399],c_w_1399);
AND_array_1506 AND_array_1506_i1400(a,b[1400],c_w_1400);
AND_array_1506 AND_array_1506_i1401(a,b[1401],c_w_1401);
AND_array_1506 AND_array_1506_i1402(a,b[1402],c_w_1402);
AND_array_1506 AND_array_1506_i1403(a,b[1403],c_w_1403);
AND_array_1506 AND_array_1506_i1404(a,b[1404],c_w_1404);
AND_array_1506 AND_array_1506_i1405(a,b[1405],c_w_1405);
AND_array_1506 AND_array_1506_i1406(a,b[1406],c_w_1406);
AND_array_1506 AND_array_1506_i1407(a,b[1407],c_w_1407);
AND_array_1506 AND_array_1506_i1408(a,b[1408],c_w_1408);
AND_array_1506 AND_array_1506_i1409(a,b[1409],c_w_1409);
AND_array_1506 AND_array_1506_i1410(a,b[1410],c_w_1410);
AND_array_1506 AND_array_1506_i1411(a,b[1411],c_w_1411);
AND_array_1506 AND_array_1506_i1412(a,b[1412],c_w_1412);
AND_array_1506 AND_array_1506_i1413(a,b[1413],c_w_1413);
AND_array_1506 AND_array_1506_i1414(a,b[1414],c_w_1414);
AND_array_1506 AND_array_1506_i1415(a,b[1415],c_w_1415);
AND_array_1506 AND_array_1506_i1416(a,b[1416],c_w_1416);
AND_array_1506 AND_array_1506_i1417(a,b[1417],c_w_1417);
AND_array_1506 AND_array_1506_i1418(a,b[1418],c_w_1418);
AND_array_1506 AND_array_1506_i1419(a,b[1419],c_w_1419);
AND_array_1506 AND_array_1506_i1420(a,b[1420],c_w_1420);
AND_array_1506 AND_array_1506_i1421(a,b[1421],c_w_1421);
AND_array_1506 AND_array_1506_i1422(a,b[1422],c_w_1422);
AND_array_1506 AND_array_1506_i1423(a,b[1423],c_w_1423);
AND_array_1506 AND_array_1506_i1424(a,b[1424],c_w_1424);
AND_array_1506 AND_array_1506_i1425(a,b[1425],c_w_1425);
AND_array_1506 AND_array_1506_i1426(a,b[1426],c_w_1426);
AND_array_1506 AND_array_1506_i1427(a,b[1427],c_w_1427);
AND_array_1506 AND_array_1506_i1428(a,b[1428],c_w_1428);
AND_array_1506 AND_array_1506_i1429(a,b[1429],c_w_1429);
AND_array_1506 AND_array_1506_i1430(a,b[1430],c_w_1430);
AND_array_1506 AND_array_1506_i1431(a,b[1431],c_w_1431);
AND_array_1506 AND_array_1506_i1432(a,b[1432],c_w_1432);
AND_array_1506 AND_array_1506_i1433(a,b[1433],c_w_1433);
AND_array_1506 AND_array_1506_i1434(a,b[1434],c_w_1434);
AND_array_1506 AND_array_1506_i1435(a,b[1435],c_w_1435);
AND_array_1506 AND_array_1506_i1436(a,b[1436],c_w_1436);
AND_array_1506 AND_array_1506_i1437(a,b[1437],c_w_1437);
AND_array_1506 AND_array_1506_i1438(a,b[1438],c_w_1438);
AND_array_1506 AND_array_1506_i1439(a,b[1439],c_w_1439);
AND_array_1506 AND_array_1506_i1440(a,b[1440],c_w_1440);
AND_array_1506 AND_array_1506_i1441(a,b[1441],c_w_1441);
AND_array_1506 AND_array_1506_i1442(a,b[1442],c_w_1442);
AND_array_1506 AND_array_1506_i1443(a,b[1443],c_w_1443);
AND_array_1506 AND_array_1506_i1444(a,b[1444],c_w_1444);
AND_array_1506 AND_array_1506_i1445(a,b[1445],c_w_1445);
AND_array_1506 AND_array_1506_i1446(a,b[1446],c_w_1446);
AND_array_1506 AND_array_1506_i1447(a,b[1447],c_w_1447);
AND_array_1506 AND_array_1506_i1448(a,b[1448],c_w_1448);
AND_array_1506 AND_array_1506_i1449(a,b[1449],c_w_1449);
AND_array_1506 AND_array_1506_i1450(a,b[1450],c_w_1450);
AND_array_1506 AND_array_1506_i1451(a,b[1451],c_w_1451);
AND_array_1506 AND_array_1506_i1452(a,b[1452],c_w_1452);
AND_array_1506 AND_array_1506_i1453(a,b[1453],c_w_1453);
AND_array_1506 AND_array_1506_i1454(a,b[1454],c_w_1454);
AND_array_1506 AND_array_1506_i1455(a,b[1455],c_w_1455);
AND_array_1506 AND_array_1506_i1456(a,b[1456],c_w_1456);
AND_array_1506 AND_array_1506_i1457(a,b[1457],c_w_1457);
AND_array_1506 AND_array_1506_i1458(a,b[1458],c_w_1458);
AND_array_1506 AND_array_1506_i1459(a,b[1459],c_w_1459);
AND_array_1506 AND_array_1506_i1460(a,b[1460],c_w_1460);
AND_array_1506 AND_array_1506_i1461(a,b[1461],c_w_1461);
AND_array_1506 AND_array_1506_i1462(a,b[1462],c_w_1462);
AND_array_1506 AND_array_1506_i1463(a,b[1463],c_w_1463);
AND_array_1506 AND_array_1506_i1464(a,b[1464],c_w_1464);
AND_array_1506 AND_array_1506_i1465(a,b[1465],c_w_1465);
AND_array_1506 AND_array_1506_i1466(a,b[1466],c_w_1466);
AND_array_1506 AND_array_1506_i1467(a,b[1467],c_w_1467);
AND_array_1506 AND_array_1506_i1468(a,b[1468],c_w_1468);
AND_array_1506 AND_array_1506_i1469(a,b[1469],c_w_1469);
AND_array_1506 AND_array_1506_i1470(a,b[1470],c_w_1470);
AND_array_1506 AND_array_1506_i1471(a,b[1471],c_w_1471);
AND_array_1506 AND_array_1506_i1472(a,b[1472],c_w_1472);
AND_array_1506 AND_array_1506_i1473(a,b[1473],c_w_1473);
AND_array_1506 AND_array_1506_i1474(a,b[1474],c_w_1474);
AND_array_1506 AND_array_1506_i1475(a,b[1475],c_w_1475);
AND_array_1506 AND_array_1506_i1476(a,b[1476],c_w_1476);
AND_array_1506 AND_array_1506_i1477(a,b[1477],c_w_1477);
AND_array_1506 AND_array_1506_i1478(a,b[1478],c_w_1478);
AND_array_1506 AND_array_1506_i1479(a,b[1479],c_w_1479);
AND_array_1506 AND_array_1506_i1480(a,b[1480],c_w_1480);
AND_array_1506 AND_array_1506_i1481(a,b[1481],c_w_1481);
AND_array_1506 AND_array_1506_i1482(a,b[1482],c_w_1482);
AND_array_1506 AND_array_1506_i1483(a,b[1483],c_w_1483);
AND_array_1506 AND_array_1506_i1484(a,b[1484],c_w_1484);
AND_array_1506 AND_array_1506_i1485(a,b[1485],c_w_1485);
AND_array_1506 AND_array_1506_i1486(a,b[1486],c_w_1486);
AND_array_1506 AND_array_1506_i1487(a,b[1487],c_w_1487);
AND_array_1506 AND_array_1506_i1488(a,b[1488],c_w_1488);
AND_array_1506 AND_array_1506_i1489(a,b[1489],c_w_1489);
AND_array_1506 AND_array_1506_i1490(a,b[1490],c_w_1490);
AND_array_1506 AND_array_1506_i1491(a,b[1491],c_w_1491);
AND_array_1506 AND_array_1506_i1492(a,b[1492],c_w_1492);
AND_array_1506 AND_array_1506_i1493(a,b[1493],c_w_1493);
AND_array_1506 AND_array_1506_i1494(a,b[1494],c_w_1494);
AND_array_1506 AND_array_1506_i1495(a,b[1495],c_w_1495);
AND_array_1506 AND_array_1506_i1496(a,b[1496],c_w_1496);
AND_array_1506 AND_array_1506_i1497(a,b[1497],c_w_1497);
AND_array_1506 AND_array_1506_i1498(a,b[1498],c_w_1498);
AND_array_1506 AND_array_1506_i1499(a,b[1499],c_w_1499);
AND_array_1506 AND_array_1506_i1500(a,b[1500],c_w_1500);
AND_array_1506 AND_array_1506_i1501(a,b[1501],c_w_1501);
AND_array_1506 AND_array_1506_i1502(a,b[1502],c_w_1502);
AND_array_1506 AND_array_1506_i1503(a,b[1503],c_w_1503);
AND_array_1506 AND_array_1506_i1504(a,b[1504],c_w_1504);
AND_array_1506 AND_array_1506_i1505(a,b[1505],c_w_1505);
    
assign c[3011:0] = {1506'b0,c_w_0};
assign c[6023:3012] = {1505'b0,c_w_1,1'b0};
assign c[9035:6024] = {1504'b0,c_w_2,2'b0};
assign c[12047:9036] = {1503'b0,c_w_3,3'b0};
assign c[15059:12048] = {1502'b0,c_w_4,4'b0};
assign c[18071:15060] = {1501'b0,c_w_5,5'b0};
assign c[21083:18072] = {1500'b0,c_w_6,6'b0};
assign c[24095:21084] = {1499'b0,c_w_7,7'b0};
assign c[27107:24096] = {1498'b0,c_w_8,8'b0};
assign c[30119:27108] = {1497'b0,c_w_9,9'b0};
assign c[33131:30120] = {1496'b0,c_w_10,10'b0};
assign c[36143:33132] = {1495'b0,c_w_11,11'b0};
assign c[39155:36144] = {1494'b0,c_w_12,12'b0};
assign c[42167:39156] = {1493'b0,c_w_13,13'b0};
assign c[45179:42168] = {1492'b0,c_w_14,14'b0};
assign c[48191:45180] = {1491'b0,c_w_15,15'b0};
assign c[51203:48192] = {1490'b0,c_w_16,16'b0};
assign c[54215:51204] = {1489'b0,c_w_17,17'b0};
assign c[57227:54216] = {1488'b0,c_w_18,18'b0};
assign c[60239:57228] = {1487'b0,c_w_19,19'b0};
assign c[63251:60240] = {1486'b0,c_w_20,20'b0};
assign c[66263:63252] = {1485'b0,c_w_21,21'b0};
assign c[69275:66264] = {1484'b0,c_w_22,22'b0};
assign c[72287:69276] = {1483'b0,c_w_23,23'b0};
assign c[75299:72288] = {1482'b0,c_w_24,24'b0};
assign c[78311:75300] = {1481'b0,c_w_25,25'b0};
assign c[81323:78312] = {1480'b0,c_w_26,26'b0};
assign c[84335:81324] = {1479'b0,c_w_27,27'b0};
assign c[87347:84336] = {1478'b0,c_w_28,28'b0};
assign c[90359:87348] = {1477'b0,c_w_29,29'b0};
assign c[93371:90360] = {1476'b0,c_w_30,30'b0};
assign c[96383:93372] = {1475'b0,c_w_31,31'b0};
assign c[99395:96384] = {1474'b0,c_w_32,32'b0};
assign c[102407:99396] = {1473'b0,c_w_33,33'b0};
assign c[105419:102408] = {1472'b0,c_w_34,34'b0};
assign c[108431:105420] = {1471'b0,c_w_35,35'b0};
assign c[111443:108432] = {1470'b0,c_w_36,36'b0};
assign c[114455:111444] = {1469'b0,c_w_37,37'b0};
assign c[117467:114456] = {1468'b0,c_w_38,38'b0};
assign c[120479:117468] = {1467'b0,c_w_39,39'b0};
assign c[123491:120480] = {1466'b0,c_w_40,40'b0};
assign c[126503:123492] = {1465'b0,c_w_41,41'b0};
assign c[129515:126504] = {1464'b0,c_w_42,42'b0};
assign c[132527:129516] = {1463'b0,c_w_43,43'b0};
assign c[135539:132528] = {1462'b0,c_w_44,44'b0};
assign c[138551:135540] = {1461'b0,c_w_45,45'b0};
assign c[141563:138552] = {1460'b0,c_w_46,46'b0};
assign c[144575:141564] = {1459'b0,c_w_47,47'b0};
assign c[147587:144576] = {1458'b0,c_w_48,48'b0};
assign c[150599:147588] = {1457'b0,c_w_49,49'b0};
assign c[153611:150600] = {1456'b0,c_w_50,50'b0};
assign c[156623:153612] = {1455'b0,c_w_51,51'b0};
assign c[159635:156624] = {1454'b0,c_w_52,52'b0};
assign c[162647:159636] = {1453'b0,c_w_53,53'b0};
assign c[165659:162648] = {1452'b0,c_w_54,54'b0};
assign c[168671:165660] = {1451'b0,c_w_55,55'b0};
assign c[171683:168672] = {1450'b0,c_w_56,56'b0};
assign c[174695:171684] = {1449'b0,c_w_57,57'b0};
assign c[177707:174696] = {1448'b0,c_w_58,58'b0};
assign c[180719:177708] = {1447'b0,c_w_59,59'b0};
assign c[183731:180720] = {1446'b0,c_w_60,60'b0};
assign c[186743:183732] = {1445'b0,c_w_61,61'b0};
assign c[189755:186744] = {1444'b0,c_w_62,62'b0};
assign c[192767:189756] = {1443'b0,c_w_63,63'b0};
assign c[195779:192768] = {1442'b0,c_w_64,64'b0};
assign c[198791:195780] = {1441'b0,c_w_65,65'b0};
assign c[201803:198792] = {1440'b0,c_w_66,66'b0};
assign c[204815:201804] = {1439'b0,c_w_67,67'b0};
assign c[207827:204816] = {1438'b0,c_w_68,68'b0};
assign c[210839:207828] = {1437'b0,c_w_69,69'b0};
assign c[213851:210840] = {1436'b0,c_w_70,70'b0};
assign c[216863:213852] = {1435'b0,c_w_71,71'b0};
assign c[219875:216864] = {1434'b0,c_w_72,72'b0};
assign c[222887:219876] = {1433'b0,c_w_73,73'b0};
assign c[225899:222888] = {1432'b0,c_w_74,74'b0};
assign c[228911:225900] = {1431'b0,c_w_75,75'b0};
assign c[231923:228912] = {1430'b0,c_w_76,76'b0};
assign c[234935:231924] = {1429'b0,c_w_77,77'b0};
assign c[237947:234936] = {1428'b0,c_w_78,78'b0};
assign c[240959:237948] = {1427'b0,c_w_79,79'b0};
assign c[243971:240960] = {1426'b0,c_w_80,80'b0};
assign c[246983:243972] = {1425'b0,c_w_81,81'b0};
assign c[249995:246984] = {1424'b0,c_w_82,82'b0};
assign c[253007:249996] = {1423'b0,c_w_83,83'b0};
assign c[256019:253008] = {1422'b0,c_w_84,84'b0};
assign c[259031:256020] = {1421'b0,c_w_85,85'b0};
assign c[262043:259032] = {1420'b0,c_w_86,86'b0};
assign c[265055:262044] = {1419'b0,c_w_87,87'b0};
assign c[268067:265056] = {1418'b0,c_w_88,88'b0};
assign c[271079:268068] = {1417'b0,c_w_89,89'b0};
assign c[274091:271080] = {1416'b0,c_w_90,90'b0};
assign c[277103:274092] = {1415'b0,c_w_91,91'b0};
assign c[280115:277104] = {1414'b0,c_w_92,92'b0};
assign c[283127:280116] = {1413'b0,c_w_93,93'b0};
assign c[286139:283128] = {1412'b0,c_w_94,94'b0};
assign c[289151:286140] = {1411'b0,c_w_95,95'b0};
assign c[292163:289152] = {1410'b0,c_w_96,96'b0};
assign c[295175:292164] = {1409'b0,c_w_97,97'b0};
assign c[298187:295176] = {1408'b0,c_w_98,98'b0};
assign c[301199:298188] = {1407'b0,c_w_99,99'b0};
assign c[304211:301200] = {1406'b0,c_w_100,100'b0};
assign c[307223:304212] = {1405'b0,c_w_101,101'b0};
assign c[310235:307224] = {1404'b0,c_w_102,102'b0};
assign c[313247:310236] = {1403'b0,c_w_103,103'b0};
assign c[316259:313248] = {1402'b0,c_w_104,104'b0};
assign c[319271:316260] = {1401'b0,c_w_105,105'b0};
assign c[322283:319272] = {1400'b0,c_w_106,106'b0};
assign c[325295:322284] = {1399'b0,c_w_107,107'b0};
assign c[328307:325296] = {1398'b0,c_w_108,108'b0};
assign c[331319:328308] = {1397'b0,c_w_109,109'b0};
assign c[334331:331320] = {1396'b0,c_w_110,110'b0};
assign c[337343:334332] = {1395'b0,c_w_111,111'b0};
assign c[340355:337344] = {1394'b0,c_w_112,112'b0};
assign c[343367:340356] = {1393'b0,c_w_113,113'b0};
assign c[346379:343368] = {1392'b0,c_w_114,114'b0};
assign c[349391:346380] = {1391'b0,c_w_115,115'b0};
assign c[352403:349392] = {1390'b0,c_w_116,116'b0};
assign c[355415:352404] = {1389'b0,c_w_117,117'b0};
assign c[358427:355416] = {1388'b0,c_w_118,118'b0};
assign c[361439:358428] = {1387'b0,c_w_119,119'b0};
assign c[364451:361440] = {1386'b0,c_w_120,120'b0};
assign c[367463:364452] = {1385'b0,c_w_121,121'b0};
assign c[370475:367464] = {1384'b0,c_w_122,122'b0};
assign c[373487:370476] = {1383'b0,c_w_123,123'b0};
assign c[376499:373488] = {1382'b0,c_w_124,124'b0};
assign c[379511:376500] = {1381'b0,c_w_125,125'b0};
assign c[382523:379512] = {1380'b0,c_w_126,126'b0};
assign c[385535:382524] = {1379'b0,c_w_127,127'b0};
assign c[388547:385536] = {1378'b0,c_w_128,128'b0};
assign c[391559:388548] = {1377'b0,c_w_129,129'b0};
assign c[394571:391560] = {1376'b0,c_w_130,130'b0};
assign c[397583:394572] = {1375'b0,c_w_131,131'b0};
assign c[400595:397584] = {1374'b0,c_w_132,132'b0};
assign c[403607:400596] = {1373'b0,c_w_133,133'b0};
assign c[406619:403608] = {1372'b0,c_w_134,134'b0};
assign c[409631:406620] = {1371'b0,c_w_135,135'b0};
assign c[412643:409632] = {1370'b0,c_w_136,136'b0};
assign c[415655:412644] = {1369'b0,c_w_137,137'b0};
assign c[418667:415656] = {1368'b0,c_w_138,138'b0};
assign c[421679:418668] = {1367'b0,c_w_139,139'b0};
assign c[424691:421680] = {1366'b0,c_w_140,140'b0};
assign c[427703:424692] = {1365'b0,c_w_141,141'b0};
assign c[430715:427704] = {1364'b0,c_w_142,142'b0};
assign c[433727:430716] = {1363'b0,c_w_143,143'b0};
assign c[436739:433728] = {1362'b0,c_w_144,144'b0};
assign c[439751:436740] = {1361'b0,c_w_145,145'b0};
assign c[442763:439752] = {1360'b0,c_w_146,146'b0};
assign c[445775:442764] = {1359'b0,c_w_147,147'b0};
assign c[448787:445776] = {1358'b0,c_w_148,148'b0};
assign c[451799:448788] = {1357'b0,c_w_149,149'b0};
assign c[454811:451800] = {1356'b0,c_w_150,150'b0};
assign c[457823:454812] = {1355'b0,c_w_151,151'b0};
assign c[460835:457824] = {1354'b0,c_w_152,152'b0};
assign c[463847:460836] = {1353'b0,c_w_153,153'b0};
assign c[466859:463848] = {1352'b0,c_w_154,154'b0};
assign c[469871:466860] = {1351'b0,c_w_155,155'b0};
assign c[472883:469872] = {1350'b0,c_w_156,156'b0};
assign c[475895:472884] = {1349'b0,c_w_157,157'b0};
assign c[478907:475896] = {1348'b0,c_w_158,158'b0};
assign c[481919:478908] = {1347'b0,c_w_159,159'b0};
assign c[484931:481920] = {1346'b0,c_w_160,160'b0};
assign c[487943:484932] = {1345'b0,c_w_161,161'b0};
assign c[490955:487944] = {1344'b0,c_w_162,162'b0};
assign c[493967:490956] = {1343'b0,c_w_163,163'b0};
assign c[496979:493968] = {1342'b0,c_w_164,164'b0};
assign c[499991:496980] = {1341'b0,c_w_165,165'b0};
assign c[503003:499992] = {1340'b0,c_w_166,166'b0};
assign c[506015:503004] = {1339'b0,c_w_167,167'b0};
assign c[509027:506016] = {1338'b0,c_w_168,168'b0};
assign c[512039:509028] = {1337'b0,c_w_169,169'b0};
assign c[515051:512040] = {1336'b0,c_w_170,170'b0};
assign c[518063:515052] = {1335'b0,c_w_171,171'b0};
assign c[521075:518064] = {1334'b0,c_w_172,172'b0};
assign c[524087:521076] = {1333'b0,c_w_173,173'b0};
assign c[527099:524088] = {1332'b0,c_w_174,174'b0};
assign c[530111:527100] = {1331'b0,c_w_175,175'b0};
assign c[533123:530112] = {1330'b0,c_w_176,176'b0};
assign c[536135:533124] = {1329'b0,c_w_177,177'b0};
assign c[539147:536136] = {1328'b0,c_w_178,178'b0};
assign c[542159:539148] = {1327'b0,c_w_179,179'b0};
assign c[545171:542160] = {1326'b0,c_w_180,180'b0};
assign c[548183:545172] = {1325'b0,c_w_181,181'b0};
assign c[551195:548184] = {1324'b0,c_w_182,182'b0};
assign c[554207:551196] = {1323'b0,c_w_183,183'b0};
assign c[557219:554208] = {1322'b0,c_w_184,184'b0};
assign c[560231:557220] = {1321'b0,c_w_185,185'b0};
assign c[563243:560232] = {1320'b0,c_w_186,186'b0};
assign c[566255:563244] = {1319'b0,c_w_187,187'b0};
assign c[569267:566256] = {1318'b0,c_w_188,188'b0};
assign c[572279:569268] = {1317'b0,c_w_189,189'b0};
assign c[575291:572280] = {1316'b0,c_w_190,190'b0};
assign c[578303:575292] = {1315'b0,c_w_191,191'b0};
assign c[581315:578304] = {1314'b0,c_w_192,192'b0};
assign c[584327:581316] = {1313'b0,c_w_193,193'b0};
assign c[587339:584328] = {1312'b0,c_w_194,194'b0};
assign c[590351:587340] = {1311'b0,c_w_195,195'b0};
assign c[593363:590352] = {1310'b0,c_w_196,196'b0};
assign c[596375:593364] = {1309'b0,c_w_197,197'b0};
assign c[599387:596376] = {1308'b0,c_w_198,198'b0};
assign c[602399:599388] = {1307'b0,c_w_199,199'b0};
assign c[605411:602400] = {1306'b0,c_w_200,200'b0};
assign c[608423:605412] = {1305'b0,c_w_201,201'b0};
assign c[611435:608424] = {1304'b0,c_w_202,202'b0};
assign c[614447:611436] = {1303'b0,c_w_203,203'b0};
assign c[617459:614448] = {1302'b0,c_w_204,204'b0};
assign c[620471:617460] = {1301'b0,c_w_205,205'b0};
assign c[623483:620472] = {1300'b0,c_w_206,206'b0};
assign c[626495:623484] = {1299'b0,c_w_207,207'b0};
assign c[629507:626496] = {1298'b0,c_w_208,208'b0};
assign c[632519:629508] = {1297'b0,c_w_209,209'b0};
assign c[635531:632520] = {1296'b0,c_w_210,210'b0};
assign c[638543:635532] = {1295'b0,c_w_211,211'b0};
assign c[641555:638544] = {1294'b0,c_w_212,212'b0};
assign c[644567:641556] = {1293'b0,c_w_213,213'b0};
assign c[647579:644568] = {1292'b0,c_w_214,214'b0};
assign c[650591:647580] = {1291'b0,c_w_215,215'b0};
assign c[653603:650592] = {1290'b0,c_w_216,216'b0};
assign c[656615:653604] = {1289'b0,c_w_217,217'b0};
assign c[659627:656616] = {1288'b0,c_w_218,218'b0};
assign c[662639:659628] = {1287'b0,c_w_219,219'b0};
assign c[665651:662640] = {1286'b0,c_w_220,220'b0};
assign c[668663:665652] = {1285'b0,c_w_221,221'b0};
assign c[671675:668664] = {1284'b0,c_w_222,222'b0};
assign c[674687:671676] = {1283'b0,c_w_223,223'b0};
assign c[677699:674688] = {1282'b0,c_w_224,224'b0};
assign c[680711:677700] = {1281'b0,c_w_225,225'b0};
assign c[683723:680712] = {1280'b0,c_w_226,226'b0};
assign c[686735:683724] = {1279'b0,c_w_227,227'b0};
assign c[689747:686736] = {1278'b0,c_w_228,228'b0};
assign c[692759:689748] = {1277'b0,c_w_229,229'b0};
assign c[695771:692760] = {1276'b0,c_w_230,230'b0};
assign c[698783:695772] = {1275'b0,c_w_231,231'b0};
assign c[701795:698784] = {1274'b0,c_w_232,232'b0};
assign c[704807:701796] = {1273'b0,c_w_233,233'b0};
assign c[707819:704808] = {1272'b0,c_w_234,234'b0};
assign c[710831:707820] = {1271'b0,c_w_235,235'b0};
assign c[713843:710832] = {1270'b0,c_w_236,236'b0};
assign c[716855:713844] = {1269'b0,c_w_237,237'b0};
assign c[719867:716856] = {1268'b0,c_w_238,238'b0};
assign c[722879:719868] = {1267'b0,c_w_239,239'b0};
assign c[725891:722880] = {1266'b0,c_w_240,240'b0};
assign c[728903:725892] = {1265'b0,c_w_241,241'b0};
assign c[731915:728904] = {1264'b0,c_w_242,242'b0};
assign c[734927:731916] = {1263'b0,c_w_243,243'b0};
assign c[737939:734928] = {1262'b0,c_w_244,244'b0};
assign c[740951:737940] = {1261'b0,c_w_245,245'b0};
assign c[743963:740952] = {1260'b0,c_w_246,246'b0};
assign c[746975:743964] = {1259'b0,c_w_247,247'b0};
assign c[749987:746976] = {1258'b0,c_w_248,248'b0};
assign c[752999:749988] = {1257'b0,c_w_249,249'b0};
assign c[756011:753000] = {1256'b0,c_w_250,250'b0};
assign c[759023:756012] = {1255'b0,c_w_251,251'b0};
assign c[762035:759024] = {1254'b0,c_w_252,252'b0};
assign c[765047:762036] = {1253'b0,c_w_253,253'b0};
assign c[768059:765048] = {1252'b0,c_w_254,254'b0};
assign c[771071:768060] = {1251'b0,c_w_255,255'b0};
assign c[774083:771072] = {1250'b0,c_w_256,256'b0};
assign c[777095:774084] = {1249'b0,c_w_257,257'b0};
assign c[780107:777096] = {1248'b0,c_w_258,258'b0};
assign c[783119:780108] = {1247'b0,c_w_259,259'b0};
assign c[786131:783120] = {1246'b0,c_w_260,260'b0};
assign c[789143:786132] = {1245'b0,c_w_261,261'b0};
assign c[792155:789144] = {1244'b0,c_w_262,262'b0};
assign c[795167:792156] = {1243'b0,c_w_263,263'b0};
assign c[798179:795168] = {1242'b0,c_w_264,264'b0};
assign c[801191:798180] = {1241'b0,c_w_265,265'b0};
assign c[804203:801192] = {1240'b0,c_w_266,266'b0};
assign c[807215:804204] = {1239'b0,c_w_267,267'b0};
assign c[810227:807216] = {1238'b0,c_w_268,268'b0};
assign c[813239:810228] = {1237'b0,c_w_269,269'b0};
assign c[816251:813240] = {1236'b0,c_w_270,270'b0};
assign c[819263:816252] = {1235'b0,c_w_271,271'b0};
assign c[822275:819264] = {1234'b0,c_w_272,272'b0};
assign c[825287:822276] = {1233'b0,c_w_273,273'b0};
assign c[828299:825288] = {1232'b0,c_w_274,274'b0};
assign c[831311:828300] = {1231'b0,c_w_275,275'b0};
assign c[834323:831312] = {1230'b0,c_w_276,276'b0};
assign c[837335:834324] = {1229'b0,c_w_277,277'b0};
assign c[840347:837336] = {1228'b0,c_w_278,278'b0};
assign c[843359:840348] = {1227'b0,c_w_279,279'b0};
assign c[846371:843360] = {1226'b0,c_w_280,280'b0};
assign c[849383:846372] = {1225'b0,c_w_281,281'b0};
assign c[852395:849384] = {1224'b0,c_w_282,282'b0};
assign c[855407:852396] = {1223'b0,c_w_283,283'b0};
assign c[858419:855408] = {1222'b0,c_w_284,284'b0};
assign c[861431:858420] = {1221'b0,c_w_285,285'b0};
assign c[864443:861432] = {1220'b0,c_w_286,286'b0};
assign c[867455:864444] = {1219'b0,c_w_287,287'b0};
assign c[870467:867456] = {1218'b0,c_w_288,288'b0};
assign c[873479:870468] = {1217'b0,c_w_289,289'b0};
assign c[876491:873480] = {1216'b0,c_w_290,290'b0};
assign c[879503:876492] = {1215'b0,c_w_291,291'b0};
assign c[882515:879504] = {1214'b0,c_w_292,292'b0};
assign c[885527:882516] = {1213'b0,c_w_293,293'b0};
assign c[888539:885528] = {1212'b0,c_w_294,294'b0};
assign c[891551:888540] = {1211'b0,c_w_295,295'b0};
assign c[894563:891552] = {1210'b0,c_w_296,296'b0};
assign c[897575:894564] = {1209'b0,c_w_297,297'b0};
assign c[900587:897576] = {1208'b0,c_w_298,298'b0};
assign c[903599:900588] = {1207'b0,c_w_299,299'b0};
assign c[906611:903600] = {1206'b0,c_w_300,300'b0};
assign c[909623:906612] = {1205'b0,c_w_301,301'b0};
assign c[912635:909624] = {1204'b0,c_w_302,302'b0};
assign c[915647:912636] = {1203'b0,c_w_303,303'b0};
assign c[918659:915648] = {1202'b0,c_w_304,304'b0};
assign c[921671:918660] = {1201'b0,c_w_305,305'b0};
assign c[924683:921672] = {1200'b0,c_w_306,306'b0};
assign c[927695:924684] = {1199'b0,c_w_307,307'b0};
assign c[930707:927696] = {1198'b0,c_w_308,308'b0};
assign c[933719:930708] = {1197'b0,c_w_309,309'b0};
assign c[936731:933720] = {1196'b0,c_w_310,310'b0};
assign c[939743:936732] = {1195'b0,c_w_311,311'b0};
assign c[942755:939744] = {1194'b0,c_w_312,312'b0};
assign c[945767:942756] = {1193'b0,c_w_313,313'b0};
assign c[948779:945768] = {1192'b0,c_w_314,314'b0};
assign c[951791:948780] = {1191'b0,c_w_315,315'b0};
assign c[954803:951792] = {1190'b0,c_w_316,316'b0};
assign c[957815:954804] = {1189'b0,c_w_317,317'b0};
assign c[960827:957816] = {1188'b0,c_w_318,318'b0};
assign c[963839:960828] = {1187'b0,c_w_319,319'b0};
assign c[966851:963840] = {1186'b0,c_w_320,320'b0};
assign c[969863:966852] = {1185'b0,c_w_321,321'b0};
assign c[972875:969864] = {1184'b0,c_w_322,322'b0};
assign c[975887:972876] = {1183'b0,c_w_323,323'b0};
assign c[978899:975888] = {1182'b0,c_w_324,324'b0};
assign c[981911:978900] = {1181'b0,c_w_325,325'b0};
assign c[984923:981912] = {1180'b0,c_w_326,326'b0};
assign c[987935:984924] = {1179'b0,c_w_327,327'b0};
assign c[990947:987936] = {1178'b0,c_w_328,328'b0};
assign c[993959:990948] = {1177'b0,c_w_329,329'b0};
assign c[996971:993960] = {1176'b0,c_w_330,330'b0};
assign c[999983:996972] = {1175'b0,c_w_331,331'b0};
assign c[1002995:999984] = {1174'b0,c_w_332,332'b0};
assign c[1006007:1002996] = {1173'b0,c_w_333,333'b0};
assign c[1009019:1006008] = {1172'b0,c_w_334,334'b0};
assign c[1012031:1009020] = {1171'b0,c_w_335,335'b0};
assign c[1015043:1012032] = {1170'b0,c_w_336,336'b0};
assign c[1018055:1015044] = {1169'b0,c_w_337,337'b0};
assign c[1021067:1018056] = {1168'b0,c_w_338,338'b0};
assign c[1024079:1021068] = {1167'b0,c_w_339,339'b0};
assign c[1027091:1024080] = {1166'b0,c_w_340,340'b0};
assign c[1030103:1027092] = {1165'b0,c_w_341,341'b0};
assign c[1033115:1030104] = {1164'b0,c_w_342,342'b0};
assign c[1036127:1033116] = {1163'b0,c_w_343,343'b0};
assign c[1039139:1036128] = {1162'b0,c_w_344,344'b0};
assign c[1042151:1039140] = {1161'b0,c_w_345,345'b0};
assign c[1045163:1042152] = {1160'b0,c_w_346,346'b0};
assign c[1048175:1045164] = {1159'b0,c_w_347,347'b0};
assign c[1051187:1048176] = {1158'b0,c_w_348,348'b0};
assign c[1054199:1051188] = {1157'b0,c_w_349,349'b0};
assign c[1057211:1054200] = {1156'b0,c_w_350,350'b0};
assign c[1060223:1057212] = {1155'b0,c_w_351,351'b0};
assign c[1063235:1060224] = {1154'b0,c_w_352,352'b0};
assign c[1066247:1063236] = {1153'b0,c_w_353,353'b0};
assign c[1069259:1066248] = {1152'b0,c_w_354,354'b0};
assign c[1072271:1069260] = {1151'b0,c_w_355,355'b0};
assign c[1075283:1072272] = {1150'b0,c_w_356,356'b0};
assign c[1078295:1075284] = {1149'b0,c_w_357,357'b0};
assign c[1081307:1078296] = {1148'b0,c_w_358,358'b0};
assign c[1084319:1081308] = {1147'b0,c_w_359,359'b0};
assign c[1087331:1084320] = {1146'b0,c_w_360,360'b0};
assign c[1090343:1087332] = {1145'b0,c_w_361,361'b0};
assign c[1093355:1090344] = {1144'b0,c_w_362,362'b0};
assign c[1096367:1093356] = {1143'b0,c_w_363,363'b0};
assign c[1099379:1096368] = {1142'b0,c_w_364,364'b0};
assign c[1102391:1099380] = {1141'b0,c_w_365,365'b0};
assign c[1105403:1102392] = {1140'b0,c_w_366,366'b0};
assign c[1108415:1105404] = {1139'b0,c_w_367,367'b0};
assign c[1111427:1108416] = {1138'b0,c_w_368,368'b0};
assign c[1114439:1111428] = {1137'b0,c_w_369,369'b0};
assign c[1117451:1114440] = {1136'b0,c_w_370,370'b0};
assign c[1120463:1117452] = {1135'b0,c_w_371,371'b0};
assign c[1123475:1120464] = {1134'b0,c_w_372,372'b0};
assign c[1126487:1123476] = {1133'b0,c_w_373,373'b0};
assign c[1129499:1126488] = {1132'b0,c_w_374,374'b0};
assign c[1132511:1129500] = {1131'b0,c_w_375,375'b0};
assign c[1135523:1132512] = {1130'b0,c_w_376,376'b0};
assign c[1138535:1135524] = {1129'b0,c_w_377,377'b0};
assign c[1141547:1138536] = {1128'b0,c_w_378,378'b0};
assign c[1144559:1141548] = {1127'b0,c_w_379,379'b0};
assign c[1147571:1144560] = {1126'b0,c_w_380,380'b0};
assign c[1150583:1147572] = {1125'b0,c_w_381,381'b0};
assign c[1153595:1150584] = {1124'b0,c_w_382,382'b0};
assign c[1156607:1153596] = {1123'b0,c_w_383,383'b0};
assign c[1159619:1156608] = {1122'b0,c_w_384,384'b0};
assign c[1162631:1159620] = {1121'b0,c_w_385,385'b0};
assign c[1165643:1162632] = {1120'b0,c_w_386,386'b0};
assign c[1168655:1165644] = {1119'b0,c_w_387,387'b0};
assign c[1171667:1168656] = {1118'b0,c_w_388,388'b0};
assign c[1174679:1171668] = {1117'b0,c_w_389,389'b0};
assign c[1177691:1174680] = {1116'b0,c_w_390,390'b0};
assign c[1180703:1177692] = {1115'b0,c_w_391,391'b0};
assign c[1183715:1180704] = {1114'b0,c_w_392,392'b0};
assign c[1186727:1183716] = {1113'b0,c_w_393,393'b0};
assign c[1189739:1186728] = {1112'b0,c_w_394,394'b0};
assign c[1192751:1189740] = {1111'b0,c_w_395,395'b0};
assign c[1195763:1192752] = {1110'b0,c_w_396,396'b0};
assign c[1198775:1195764] = {1109'b0,c_w_397,397'b0};
assign c[1201787:1198776] = {1108'b0,c_w_398,398'b0};
assign c[1204799:1201788] = {1107'b0,c_w_399,399'b0};
assign c[1207811:1204800] = {1106'b0,c_w_400,400'b0};
assign c[1210823:1207812] = {1105'b0,c_w_401,401'b0};
assign c[1213835:1210824] = {1104'b0,c_w_402,402'b0};
assign c[1216847:1213836] = {1103'b0,c_w_403,403'b0};
assign c[1219859:1216848] = {1102'b0,c_w_404,404'b0};
assign c[1222871:1219860] = {1101'b0,c_w_405,405'b0};
assign c[1225883:1222872] = {1100'b0,c_w_406,406'b0};
assign c[1228895:1225884] = {1099'b0,c_w_407,407'b0};
assign c[1231907:1228896] = {1098'b0,c_w_408,408'b0};
assign c[1234919:1231908] = {1097'b0,c_w_409,409'b0};
assign c[1237931:1234920] = {1096'b0,c_w_410,410'b0};
assign c[1240943:1237932] = {1095'b0,c_w_411,411'b0};
assign c[1243955:1240944] = {1094'b0,c_w_412,412'b0};
assign c[1246967:1243956] = {1093'b0,c_w_413,413'b0};
assign c[1249979:1246968] = {1092'b0,c_w_414,414'b0};
assign c[1252991:1249980] = {1091'b0,c_w_415,415'b0};
assign c[1256003:1252992] = {1090'b0,c_w_416,416'b0};
assign c[1259015:1256004] = {1089'b0,c_w_417,417'b0};
assign c[1262027:1259016] = {1088'b0,c_w_418,418'b0};
assign c[1265039:1262028] = {1087'b0,c_w_419,419'b0};
assign c[1268051:1265040] = {1086'b0,c_w_420,420'b0};
assign c[1271063:1268052] = {1085'b0,c_w_421,421'b0};
assign c[1274075:1271064] = {1084'b0,c_w_422,422'b0};
assign c[1277087:1274076] = {1083'b0,c_w_423,423'b0};
assign c[1280099:1277088] = {1082'b0,c_w_424,424'b0};
assign c[1283111:1280100] = {1081'b0,c_w_425,425'b0};
assign c[1286123:1283112] = {1080'b0,c_w_426,426'b0};
assign c[1289135:1286124] = {1079'b0,c_w_427,427'b0};
assign c[1292147:1289136] = {1078'b0,c_w_428,428'b0};
assign c[1295159:1292148] = {1077'b0,c_w_429,429'b0};
assign c[1298171:1295160] = {1076'b0,c_w_430,430'b0};
assign c[1301183:1298172] = {1075'b0,c_w_431,431'b0};
assign c[1304195:1301184] = {1074'b0,c_w_432,432'b0};
assign c[1307207:1304196] = {1073'b0,c_w_433,433'b0};
assign c[1310219:1307208] = {1072'b0,c_w_434,434'b0};
assign c[1313231:1310220] = {1071'b0,c_w_435,435'b0};
assign c[1316243:1313232] = {1070'b0,c_w_436,436'b0};
assign c[1319255:1316244] = {1069'b0,c_w_437,437'b0};
assign c[1322267:1319256] = {1068'b0,c_w_438,438'b0};
assign c[1325279:1322268] = {1067'b0,c_w_439,439'b0};
assign c[1328291:1325280] = {1066'b0,c_w_440,440'b0};
assign c[1331303:1328292] = {1065'b0,c_w_441,441'b0};
assign c[1334315:1331304] = {1064'b0,c_w_442,442'b0};
assign c[1337327:1334316] = {1063'b0,c_w_443,443'b0};
assign c[1340339:1337328] = {1062'b0,c_w_444,444'b0};
assign c[1343351:1340340] = {1061'b0,c_w_445,445'b0};
assign c[1346363:1343352] = {1060'b0,c_w_446,446'b0};
assign c[1349375:1346364] = {1059'b0,c_w_447,447'b0};
assign c[1352387:1349376] = {1058'b0,c_w_448,448'b0};
assign c[1355399:1352388] = {1057'b0,c_w_449,449'b0};
assign c[1358411:1355400] = {1056'b0,c_w_450,450'b0};
assign c[1361423:1358412] = {1055'b0,c_w_451,451'b0};
assign c[1364435:1361424] = {1054'b0,c_w_452,452'b0};
assign c[1367447:1364436] = {1053'b0,c_w_453,453'b0};
assign c[1370459:1367448] = {1052'b0,c_w_454,454'b0};
assign c[1373471:1370460] = {1051'b0,c_w_455,455'b0};
assign c[1376483:1373472] = {1050'b0,c_w_456,456'b0};
assign c[1379495:1376484] = {1049'b0,c_w_457,457'b0};
assign c[1382507:1379496] = {1048'b0,c_w_458,458'b0};
assign c[1385519:1382508] = {1047'b0,c_w_459,459'b0};
assign c[1388531:1385520] = {1046'b0,c_w_460,460'b0};
assign c[1391543:1388532] = {1045'b0,c_w_461,461'b0};
assign c[1394555:1391544] = {1044'b0,c_w_462,462'b0};
assign c[1397567:1394556] = {1043'b0,c_w_463,463'b0};
assign c[1400579:1397568] = {1042'b0,c_w_464,464'b0};
assign c[1403591:1400580] = {1041'b0,c_w_465,465'b0};
assign c[1406603:1403592] = {1040'b0,c_w_466,466'b0};
assign c[1409615:1406604] = {1039'b0,c_w_467,467'b0};
assign c[1412627:1409616] = {1038'b0,c_w_468,468'b0};
assign c[1415639:1412628] = {1037'b0,c_w_469,469'b0};
assign c[1418651:1415640] = {1036'b0,c_w_470,470'b0};
assign c[1421663:1418652] = {1035'b0,c_w_471,471'b0};
assign c[1424675:1421664] = {1034'b0,c_w_472,472'b0};
assign c[1427687:1424676] = {1033'b0,c_w_473,473'b0};
assign c[1430699:1427688] = {1032'b0,c_w_474,474'b0};
assign c[1433711:1430700] = {1031'b0,c_w_475,475'b0};
assign c[1436723:1433712] = {1030'b0,c_w_476,476'b0};
assign c[1439735:1436724] = {1029'b0,c_w_477,477'b0};
assign c[1442747:1439736] = {1028'b0,c_w_478,478'b0};
assign c[1445759:1442748] = {1027'b0,c_w_479,479'b0};
assign c[1448771:1445760] = {1026'b0,c_w_480,480'b0};
assign c[1451783:1448772] = {1025'b0,c_w_481,481'b0};
assign c[1454795:1451784] = {1024'b0,c_w_482,482'b0};
assign c[1457807:1454796] = {1023'b0,c_w_483,483'b0};
assign c[1460819:1457808] = {1022'b0,c_w_484,484'b0};
assign c[1463831:1460820] = {1021'b0,c_w_485,485'b0};
assign c[1466843:1463832] = {1020'b0,c_w_486,486'b0};
assign c[1469855:1466844] = {1019'b0,c_w_487,487'b0};
assign c[1472867:1469856] = {1018'b0,c_w_488,488'b0};
assign c[1475879:1472868] = {1017'b0,c_w_489,489'b0};
assign c[1478891:1475880] = {1016'b0,c_w_490,490'b0};
assign c[1481903:1478892] = {1015'b0,c_w_491,491'b0};
assign c[1484915:1481904] = {1014'b0,c_w_492,492'b0};
assign c[1487927:1484916] = {1013'b0,c_w_493,493'b0};
assign c[1490939:1487928] = {1012'b0,c_w_494,494'b0};
assign c[1493951:1490940] = {1011'b0,c_w_495,495'b0};
assign c[1496963:1493952] = {1010'b0,c_w_496,496'b0};
assign c[1499975:1496964] = {1009'b0,c_w_497,497'b0};
assign c[1502987:1499976] = {1008'b0,c_w_498,498'b0};
assign c[1505999:1502988] = {1007'b0,c_w_499,499'b0};
assign c[1509011:1506000] = {1006'b0,c_w_500,500'b0};
assign c[1512023:1509012] = {1005'b0,c_w_501,501'b0};
assign c[1515035:1512024] = {1004'b0,c_w_502,502'b0};
assign c[1518047:1515036] = {1003'b0,c_w_503,503'b0};
assign c[1521059:1518048] = {1002'b0,c_w_504,504'b0};
assign c[1524071:1521060] = {1001'b0,c_w_505,505'b0};
assign c[1527083:1524072] = {1000'b0,c_w_506,506'b0};
assign c[1530095:1527084] = {999'b0,c_w_507,507'b0};
assign c[1533107:1530096] = {998'b0,c_w_508,508'b0};
assign c[1536119:1533108] = {997'b0,c_w_509,509'b0};
assign c[1539131:1536120] = {996'b0,c_w_510,510'b0};
assign c[1542143:1539132] = {995'b0,c_w_511,511'b0};
assign c[1545155:1542144] = {994'b0,c_w_512,512'b0};
assign c[1548167:1545156] = {993'b0,c_w_513,513'b0};
assign c[1551179:1548168] = {992'b0,c_w_514,514'b0};
assign c[1554191:1551180] = {991'b0,c_w_515,515'b0};
assign c[1557203:1554192] = {990'b0,c_w_516,516'b0};
assign c[1560215:1557204] = {989'b0,c_w_517,517'b0};
assign c[1563227:1560216] = {988'b0,c_w_518,518'b0};
assign c[1566239:1563228] = {987'b0,c_w_519,519'b0};
assign c[1569251:1566240] = {986'b0,c_w_520,520'b0};
assign c[1572263:1569252] = {985'b0,c_w_521,521'b0};
assign c[1575275:1572264] = {984'b0,c_w_522,522'b0};
assign c[1578287:1575276] = {983'b0,c_w_523,523'b0};
assign c[1581299:1578288] = {982'b0,c_w_524,524'b0};
assign c[1584311:1581300] = {981'b0,c_w_525,525'b0};
assign c[1587323:1584312] = {980'b0,c_w_526,526'b0};
assign c[1590335:1587324] = {979'b0,c_w_527,527'b0};
assign c[1593347:1590336] = {978'b0,c_w_528,528'b0};
assign c[1596359:1593348] = {977'b0,c_w_529,529'b0};
assign c[1599371:1596360] = {976'b0,c_w_530,530'b0};
assign c[1602383:1599372] = {975'b0,c_w_531,531'b0};
assign c[1605395:1602384] = {974'b0,c_w_532,532'b0};
assign c[1608407:1605396] = {973'b0,c_w_533,533'b0};
assign c[1611419:1608408] = {972'b0,c_w_534,534'b0};
assign c[1614431:1611420] = {971'b0,c_w_535,535'b0};
assign c[1617443:1614432] = {970'b0,c_w_536,536'b0};
assign c[1620455:1617444] = {969'b0,c_w_537,537'b0};
assign c[1623467:1620456] = {968'b0,c_w_538,538'b0};
assign c[1626479:1623468] = {967'b0,c_w_539,539'b0};
assign c[1629491:1626480] = {966'b0,c_w_540,540'b0};
assign c[1632503:1629492] = {965'b0,c_w_541,541'b0};
assign c[1635515:1632504] = {964'b0,c_w_542,542'b0};
assign c[1638527:1635516] = {963'b0,c_w_543,543'b0};
assign c[1641539:1638528] = {962'b0,c_w_544,544'b0};
assign c[1644551:1641540] = {961'b0,c_w_545,545'b0};
assign c[1647563:1644552] = {960'b0,c_w_546,546'b0};
assign c[1650575:1647564] = {959'b0,c_w_547,547'b0};
assign c[1653587:1650576] = {958'b0,c_w_548,548'b0};
assign c[1656599:1653588] = {957'b0,c_w_549,549'b0};
assign c[1659611:1656600] = {956'b0,c_w_550,550'b0};
assign c[1662623:1659612] = {955'b0,c_w_551,551'b0};
assign c[1665635:1662624] = {954'b0,c_w_552,552'b0};
assign c[1668647:1665636] = {953'b0,c_w_553,553'b0};
assign c[1671659:1668648] = {952'b0,c_w_554,554'b0};
assign c[1674671:1671660] = {951'b0,c_w_555,555'b0};
assign c[1677683:1674672] = {950'b0,c_w_556,556'b0};
assign c[1680695:1677684] = {949'b0,c_w_557,557'b0};
assign c[1683707:1680696] = {948'b0,c_w_558,558'b0};
assign c[1686719:1683708] = {947'b0,c_w_559,559'b0};
assign c[1689731:1686720] = {946'b0,c_w_560,560'b0};
assign c[1692743:1689732] = {945'b0,c_w_561,561'b0};
assign c[1695755:1692744] = {944'b0,c_w_562,562'b0};
assign c[1698767:1695756] = {943'b0,c_w_563,563'b0};
assign c[1701779:1698768] = {942'b0,c_w_564,564'b0};
assign c[1704791:1701780] = {941'b0,c_w_565,565'b0};
assign c[1707803:1704792] = {940'b0,c_w_566,566'b0};
assign c[1710815:1707804] = {939'b0,c_w_567,567'b0};
assign c[1713827:1710816] = {938'b0,c_w_568,568'b0};
assign c[1716839:1713828] = {937'b0,c_w_569,569'b0};
assign c[1719851:1716840] = {936'b0,c_w_570,570'b0};
assign c[1722863:1719852] = {935'b0,c_w_571,571'b0};
assign c[1725875:1722864] = {934'b0,c_w_572,572'b0};
assign c[1728887:1725876] = {933'b0,c_w_573,573'b0};
assign c[1731899:1728888] = {932'b0,c_w_574,574'b0};
assign c[1734911:1731900] = {931'b0,c_w_575,575'b0};
assign c[1737923:1734912] = {930'b0,c_w_576,576'b0};
assign c[1740935:1737924] = {929'b0,c_w_577,577'b0};
assign c[1743947:1740936] = {928'b0,c_w_578,578'b0};
assign c[1746959:1743948] = {927'b0,c_w_579,579'b0};
assign c[1749971:1746960] = {926'b0,c_w_580,580'b0};
assign c[1752983:1749972] = {925'b0,c_w_581,581'b0};
assign c[1755995:1752984] = {924'b0,c_w_582,582'b0};
assign c[1759007:1755996] = {923'b0,c_w_583,583'b0};
assign c[1762019:1759008] = {922'b0,c_w_584,584'b0};
assign c[1765031:1762020] = {921'b0,c_w_585,585'b0};
assign c[1768043:1765032] = {920'b0,c_w_586,586'b0};
assign c[1771055:1768044] = {919'b0,c_w_587,587'b0};
assign c[1774067:1771056] = {918'b0,c_w_588,588'b0};
assign c[1777079:1774068] = {917'b0,c_w_589,589'b0};
assign c[1780091:1777080] = {916'b0,c_w_590,590'b0};
assign c[1783103:1780092] = {915'b0,c_w_591,591'b0};
assign c[1786115:1783104] = {914'b0,c_w_592,592'b0};
assign c[1789127:1786116] = {913'b0,c_w_593,593'b0};
assign c[1792139:1789128] = {912'b0,c_w_594,594'b0};
assign c[1795151:1792140] = {911'b0,c_w_595,595'b0};
assign c[1798163:1795152] = {910'b0,c_w_596,596'b0};
assign c[1801175:1798164] = {909'b0,c_w_597,597'b0};
assign c[1804187:1801176] = {908'b0,c_w_598,598'b0};
assign c[1807199:1804188] = {907'b0,c_w_599,599'b0};
assign c[1810211:1807200] = {906'b0,c_w_600,600'b0};
assign c[1813223:1810212] = {905'b0,c_w_601,601'b0};
assign c[1816235:1813224] = {904'b0,c_w_602,602'b0};
assign c[1819247:1816236] = {903'b0,c_w_603,603'b0};
assign c[1822259:1819248] = {902'b0,c_w_604,604'b0};
assign c[1825271:1822260] = {901'b0,c_w_605,605'b0};
assign c[1828283:1825272] = {900'b0,c_w_606,606'b0};
assign c[1831295:1828284] = {899'b0,c_w_607,607'b0};
assign c[1834307:1831296] = {898'b0,c_w_608,608'b0};
assign c[1837319:1834308] = {897'b0,c_w_609,609'b0};
assign c[1840331:1837320] = {896'b0,c_w_610,610'b0};
assign c[1843343:1840332] = {895'b0,c_w_611,611'b0};
assign c[1846355:1843344] = {894'b0,c_w_612,612'b0};
assign c[1849367:1846356] = {893'b0,c_w_613,613'b0};
assign c[1852379:1849368] = {892'b0,c_w_614,614'b0};
assign c[1855391:1852380] = {891'b0,c_w_615,615'b0};
assign c[1858403:1855392] = {890'b0,c_w_616,616'b0};
assign c[1861415:1858404] = {889'b0,c_w_617,617'b0};
assign c[1864427:1861416] = {888'b0,c_w_618,618'b0};
assign c[1867439:1864428] = {887'b0,c_w_619,619'b0};
assign c[1870451:1867440] = {886'b0,c_w_620,620'b0};
assign c[1873463:1870452] = {885'b0,c_w_621,621'b0};
assign c[1876475:1873464] = {884'b0,c_w_622,622'b0};
assign c[1879487:1876476] = {883'b0,c_w_623,623'b0};
assign c[1882499:1879488] = {882'b0,c_w_624,624'b0};
assign c[1885511:1882500] = {881'b0,c_w_625,625'b0};
assign c[1888523:1885512] = {880'b0,c_w_626,626'b0};
assign c[1891535:1888524] = {879'b0,c_w_627,627'b0};
assign c[1894547:1891536] = {878'b0,c_w_628,628'b0};
assign c[1897559:1894548] = {877'b0,c_w_629,629'b0};
assign c[1900571:1897560] = {876'b0,c_w_630,630'b0};
assign c[1903583:1900572] = {875'b0,c_w_631,631'b0};
assign c[1906595:1903584] = {874'b0,c_w_632,632'b0};
assign c[1909607:1906596] = {873'b0,c_w_633,633'b0};
assign c[1912619:1909608] = {872'b0,c_w_634,634'b0};
assign c[1915631:1912620] = {871'b0,c_w_635,635'b0};
assign c[1918643:1915632] = {870'b0,c_w_636,636'b0};
assign c[1921655:1918644] = {869'b0,c_w_637,637'b0};
assign c[1924667:1921656] = {868'b0,c_w_638,638'b0};
assign c[1927679:1924668] = {867'b0,c_w_639,639'b0};
assign c[1930691:1927680] = {866'b0,c_w_640,640'b0};
assign c[1933703:1930692] = {865'b0,c_w_641,641'b0};
assign c[1936715:1933704] = {864'b0,c_w_642,642'b0};
assign c[1939727:1936716] = {863'b0,c_w_643,643'b0};
assign c[1942739:1939728] = {862'b0,c_w_644,644'b0};
assign c[1945751:1942740] = {861'b0,c_w_645,645'b0};
assign c[1948763:1945752] = {860'b0,c_w_646,646'b0};
assign c[1951775:1948764] = {859'b0,c_w_647,647'b0};
assign c[1954787:1951776] = {858'b0,c_w_648,648'b0};
assign c[1957799:1954788] = {857'b0,c_w_649,649'b0};
assign c[1960811:1957800] = {856'b0,c_w_650,650'b0};
assign c[1963823:1960812] = {855'b0,c_w_651,651'b0};
assign c[1966835:1963824] = {854'b0,c_w_652,652'b0};
assign c[1969847:1966836] = {853'b0,c_w_653,653'b0};
assign c[1972859:1969848] = {852'b0,c_w_654,654'b0};
assign c[1975871:1972860] = {851'b0,c_w_655,655'b0};
assign c[1978883:1975872] = {850'b0,c_w_656,656'b0};
assign c[1981895:1978884] = {849'b0,c_w_657,657'b0};
assign c[1984907:1981896] = {848'b0,c_w_658,658'b0};
assign c[1987919:1984908] = {847'b0,c_w_659,659'b0};
assign c[1990931:1987920] = {846'b0,c_w_660,660'b0};
assign c[1993943:1990932] = {845'b0,c_w_661,661'b0};
assign c[1996955:1993944] = {844'b0,c_w_662,662'b0};
assign c[1999967:1996956] = {843'b0,c_w_663,663'b0};
assign c[2002979:1999968] = {842'b0,c_w_664,664'b0};
assign c[2005991:2002980] = {841'b0,c_w_665,665'b0};
assign c[2009003:2005992] = {840'b0,c_w_666,666'b0};
assign c[2012015:2009004] = {839'b0,c_w_667,667'b0};
assign c[2015027:2012016] = {838'b0,c_w_668,668'b0};
assign c[2018039:2015028] = {837'b0,c_w_669,669'b0};
assign c[2021051:2018040] = {836'b0,c_w_670,670'b0};
assign c[2024063:2021052] = {835'b0,c_w_671,671'b0};
assign c[2027075:2024064] = {834'b0,c_w_672,672'b0};
assign c[2030087:2027076] = {833'b0,c_w_673,673'b0};
assign c[2033099:2030088] = {832'b0,c_w_674,674'b0};
assign c[2036111:2033100] = {831'b0,c_w_675,675'b0};
assign c[2039123:2036112] = {830'b0,c_w_676,676'b0};
assign c[2042135:2039124] = {829'b0,c_w_677,677'b0};
assign c[2045147:2042136] = {828'b0,c_w_678,678'b0};
assign c[2048159:2045148] = {827'b0,c_w_679,679'b0};
assign c[2051171:2048160] = {826'b0,c_w_680,680'b0};
assign c[2054183:2051172] = {825'b0,c_w_681,681'b0};
assign c[2057195:2054184] = {824'b0,c_w_682,682'b0};
assign c[2060207:2057196] = {823'b0,c_w_683,683'b0};
assign c[2063219:2060208] = {822'b0,c_w_684,684'b0};
assign c[2066231:2063220] = {821'b0,c_w_685,685'b0};
assign c[2069243:2066232] = {820'b0,c_w_686,686'b0};
assign c[2072255:2069244] = {819'b0,c_w_687,687'b0};
assign c[2075267:2072256] = {818'b0,c_w_688,688'b0};
assign c[2078279:2075268] = {817'b0,c_w_689,689'b0};
assign c[2081291:2078280] = {816'b0,c_w_690,690'b0};
assign c[2084303:2081292] = {815'b0,c_w_691,691'b0};
assign c[2087315:2084304] = {814'b0,c_w_692,692'b0};
assign c[2090327:2087316] = {813'b0,c_w_693,693'b0};
assign c[2093339:2090328] = {812'b0,c_w_694,694'b0};
assign c[2096351:2093340] = {811'b0,c_w_695,695'b0};
assign c[2099363:2096352] = {810'b0,c_w_696,696'b0};
assign c[2102375:2099364] = {809'b0,c_w_697,697'b0};
assign c[2105387:2102376] = {808'b0,c_w_698,698'b0};
assign c[2108399:2105388] = {807'b0,c_w_699,699'b0};
assign c[2111411:2108400] = {806'b0,c_w_700,700'b0};
assign c[2114423:2111412] = {805'b0,c_w_701,701'b0};
assign c[2117435:2114424] = {804'b0,c_w_702,702'b0};
assign c[2120447:2117436] = {803'b0,c_w_703,703'b0};
assign c[2123459:2120448] = {802'b0,c_w_704,704'b0};
assign c[2126471:2123460] = {801'b0,c_w_705,705'b0};
assign c[2129483:2126472] = {800'b0,c_w_706,706'b0};
assign c[2132495:2129484] = {799'b0,c_w_707,707'b0};
assign c[2135507:2132496] = {798'b0,c_w_708,708'b0};
assign c[2138519:2135508] = {797'b0,c_w_709,709'b0};
assign c[2141531:2138520] = {796'b0,c_w_710,710'b0};
assign c[2144543:2141532] = {795'b0,c_w_711,711'b0};
assign c[2147555:2144544] = {794'b0,c_w_712,712'b0};
assign c[2150567:2147556] = {793'b0,c_w_713,713'b0};
assign c[2153579:2150568] = {792'b0,c_w_714,714'b0};
assign c[2156591:2153580] = {791'b0,c_w_715,715'b0};
assign c[2159603:2156592] = {790'b0,c_w_716,716'b0};
assign c[2162615:2159604] = {789'b0,c_w_717,717'b0};
assign c[2165627:2162616] = {788'b0,c_w_718,718'b0};
assign c[2168639:2165628] = {787'b0,c_w_719,719'b0};
assign c[2171651:2168640] = {786'b0,c_w_720,720'b0};
assign c[2174663:2171652] = {785'b0,c_w_721,721'b0};
assign c[2177675:2174664] = {784'b0,c_w_722,722'b0};
assign c[2180687:2177676] = {783'b0,c_w_723,723'b0};
assign c[2183699:2180688] = {782'b0,c_w_724,724'b0};
assign c[2186711:2183700] = {781'b0,c_w_725,725'b0};
assign c[2189723:2186712] = {780'b0,c_w_726,726'b0};
assign c[2192735:2189724] = {779'b0,c_w_727,727'b0};
assign c[2195747:2192736] = {778'b0,c_w_728,728'b0};
assign c[2198759:2195748] = {777'b0,c_w_729,729'b0};
assign c[2201771:2198760] = {776'b0,c_w_730,730'b0};
assign c[2204783:2201772] = {775'b0,c_w_731,731'b0};
assign c[2207795:2204784] = {774'b0,c_w_732,732'b0};
assign c[2210807:2207796] = {773'b0,c_w_733,733'b0};
assign c[2213819:2210808] = {772'b0,c_w_734,734'b0};
assign c[2216831:2213820] = {771'b0,c_w_735,735'b0};
assign c[2219843:2216832] = {770'b0,c_w_736,736'b0};
assign c[2222855:2219844] = {769'b0,c_w_737,737'b0};
assign c[2225867:2222856] = {768'b0,c_w_738,738'b0};
assign c[2228879:2225868] = {767'b0,c_w_739,739'b0};
assign c[2231891:2228880] = {766'b0,c_w_740,740'b0};
assign c[2234903:2231892] = {765'b0,c_w_741,741'b0};
assign c[2237915:2234904] = {764'b0,c_w_742,742'b0};
assign c[2240927:2237916] = {763'b0,c_w_743,743'b0};
assign c[2243939:2240928] = {762'b0,c_w_744,744'b0};
assign c[2246951:2243940] = {761'b0,c_w_745,745'b0};
assign c[2249963:2246952] = {760'b0,c_w_746,746'b0};
assign c[2252975:2249964] = {759'b0,c_w_747,747'b0};
assign c[2255987:2252976] = {758'b0,c_w_748,748'b0};
assign c[2258999:2255988] = {757'b0,c_w_749,749'b0};
assign c[2262011:2259000] = {756'b0,c_w_750,750'b0};
assign c[2265023:2262012] = {755'b0,c_w_751,751'b0};
assign c[2268035:2265024] = {754'b0,c_w_752,752'b0};
assign c[2271047:2268036] = {753'b0,c_w_753,753'b0};
assign c[2274059:2271048] = {752'b0,c_w_754,754'b0};
assign c[2277071:2274060] = {751'b0,c_w_755,755'b0};
assign c[2280083:2277072] = {750'b0,c_w_756,756'b0};
assign c[2283095:2280084] = {749'b0,c_w_757,757'b0};
assign c[2286107:2283096] = {748'b0,c_w_758,758'b0};
assign c[2289119:2286108] = {747'b0,c_w_759,759'b0};
assign c[2292131:2289120] = {746'b0,c_w_760,760'b0};
assign c[2295143:2292132] = {745'b0,c_w_761,761'b0};
assign c[2298155:2295144] = {744'b0,c_w_762,762'b0};
assign c[2301167:2298156] = {743'b0,c_w_763,763'b0};
assign c[2304179:2301168] = {742'b0,c_w_764,764'b0};
assign c[2307191:2304180] = {741'b0,c_w_765,765'b0};
assign c[2310203:2307192] = {740'b0,c_w_766,766'b0};
assign c[2313215:2310204] = {739'b0,c_w_767,767'b0};
assign c[2316227:2313216] = {738'b0,c_w_768,768'b0};
assign c[2319239:2316228] = {737'b0,c_w_769,769'b0};
assign c[2322251:2319240] = {736'b0,c_w_770,770'b0};
assign c[2325263:2322252] = {735'b0,c_w_771,771'b0};
assign c[2328275:2325264] = {734'b0,c_w_772,772'b0};
assign c[2331287:2328276] = {733'b0,c_w_773,773'b0};
assign c[2334299:2331288] = {732'b0,c_w_774,774'b0};
assign c[2337311:2334300] = {731'b0,c_w_775,775'b0};
assign c[2340323:2337312] = {730'b0,c_w_776,776'b0};
assign c[2343335:2340324] = {729'b0,c_w_777,777'b0};
assign c[2346347:2343336] = {728'b0,c_w_778,778'b0};
assign c[2349359:2346348] = {727'b0,c_w_779,779'b0};
assign c[2352371:2349360] = {726'b0,c_w_780,780'b0};
assign c[2355383:2352372] = {725'b0,c_w_781,781'b0};
assign c[2358395:2355384] = {724'b0,c_w_782,782'b0};
assign c[2361407:2358396] = {723'b0,c_w_783,783'b0};
assign c[2364419:2361408] = {722'b0,c_w_784,784'b0};
assign c[2367431:2364420] = {721'b0,c_w_785,785'b0};
assign c[2370443:2367432] = {720'b0,c_w_786,786'b0};
assign c[2373455:2370444] = {719'b0,c_w_787,787'b0};
assign c[2376467:2373456] = {718'b0,c_w_788,788'b0};
assign c[2379479:2376468] = {717'b0,c_w_789,789'b0};
assign c[2382491:2379480] = {716'b0,c_w_790,790'b0};
assign c[2385503:2382492] = {715'b0,c_w_791,791'b0};
assign c[2388515:2385504] = {714'b0,c_w_792,792'b0};
assign c[2391527:2388516] = {713'b0,c_w_793,793'b0};
assign c[2394539:2391528] = {712'b0,c_w_794,794'b0};
assign c[2397551:2394540] = {711'b0,c_w_795,795'b0};
assign c[2400563:2397552] = {710'b0,c_w_796,796'b0};
assign c[2403575:2400564] = {709'b0,c_w_797,797'b0};
assign c[2406587:2403576] = {708'b0,c_w_798,798'b0};
assign c[2409599:2406588] = {707'b0,c_w_799,799'b0};
assign c[2412611:2409600] = {706'b0,c_w_800,800'b0};
assign c[2415623:2412612] = {705'b0,c_w_801,801'b0};
assign c[2418635:2415624] = {704'b0,c_w_802,802'b0};
assign c[2421647:2418636] = {703'b0,c_w_803,803'b0};
assign c[2424659:2421648] = {702'b0,c_w_804,804'b0};
assign c[2427671:2424660] = {701'b0,c_w_805,805'b0};
assign c[2430683:2427672] = {700'b0,c_w_806,806'b0};
assign c[2433695:2430684] = {699'b0,c_w_807,807'b0};
assign c[2436707:2433696] = {698'b0,c_w_808,808'b0};
assign c[2439719:2436708] = {697'b0,c_w_809,809'b0};
assign c[2442731:2439720] = {696'b0,c_w_810,810'b0};
assign c[2445743:2442732] = {695'b0,c_w_811,811'b0};
assign c[2448755:2445744] = {694'b0,c_w_812,812'b0};
assign c[2451767:2448756] = {693'b0,c_w_813,813'b0};
assign c[2454779:2451768] = {692'b0,c_w_814,814'b0};
assign c[2457791:2454780] = {691'b0,c_w_815,815'b0};
assign c[2460803:2457792] = {690'b0,c_w_816,816'b0};
assign c[2463815:2460804] = {689'b0,c_w_817,817'b0};
assign c[2466827:2463816] = {688'b0,c_w_818,818'b0};
assign c[2469839:2466828] = {687'b0,c_w_819,819'b0};
assign c[2472851:2469840] = {686'b0,c_w_820,820'b0};
assign c[2475863:2472852] = {685'b0,c_w_821,821'b0};
assign c[2478875:2475864] = {684'b0,c_w_822,822'b0};
assign c[2481887:2478876] = {683'b0,c_w_823,823'b0};
assign c[2484899:2481888] = {682'b0,c_w_824,824'b0};
assign c[2487911:2484900] = {681'b0,c_w_825,825'b0};
assign c[2490923:2487912] = {680'b0,c_w_826,826'b0};
assign c[2493935:2490924] = {679'b0,c_w_827,827'b0};
assign c[2496947:2493936] = {678'b0,c_w_828,828'b0};
assign c[2499959:2496948] = {677'b0,c_w_829,829'b0};
assign c[2502971:2499960] = {676'b0,c_w_830,830'b0};
assign c[2505983:2502972] = {675'b0,c_w_831,831'b0};
assign c[2508995:2505984] = {674'b0,c_w_832,832'b0};
assign c[2512007:2508996] = {673'b0,c_w_833,833'b0};
assign c[2515019:2512008] = {672'b0,c_w_834,834'b0};
assign c[2518031:2515020] = {671'b0,c_w_835,835'b0};
assign c[2521043:2518032] = {670'b0,c_w_836,836'b0};
assign c[2524055:2521044] = {669'b0,c_w_837,837'b0};
assign c[2527067:2524056] = {668'b0,c_w_838,838'b0};
assign c[2530079:2527068] = {667'b0,c_w_839,839'b0};
assign c[2533091:2530080] = {666'b0,c_w_840,840'b0};
assign c[2536103:2533092] = {665'b0,c_w_841,841'b0};
assign c[2539115:2536104] = {664'b0,c_w_842,842'b0};
assign c[2542127:2539116] = {663'b0,c_w_843,843'b0};
assign c[2545139:2542128] = {662'b0,c_w_844,844'b0};
assign c[2548151:2545140] = {661'b0,c_w_845,845'b0};
assign c[2551163:2548152] = {660'b0,c_w_846,846'b0};
assign c[2554175:2551164] = {659'b0,c_w_847,847'b0};
assign c[2557187:2554176] = {658'b0,c_w_848,848'b0};
assign c[2560199:2557188] = {657'b0,c_w_849,849'b0};
assign c[2563211:2560200] = {656'b0,c_w_850,850'b0};
assign c[2566223:2563212] = {655'b0,c_w_851,851'b0};
assign c[2569235:2566224] = {654'b0,c_w_852,852'b0};
assign c[2572247:2569236] = {653'b0,c_w_853,853'b0};
assign c[2575259:2572248] = {652'b0,c_w_854,854'b0};
assign c[2578271:2575260] = {651'b0,c_w_855,855'b0};
assign c[2581283:2578272] = {650'b0,c_w_856,856'b0};
assign c[2584295:2581284] = {649'b0,c_w_857,857'b0};
assign c[2587307:2584296] = {648'b0,c_w_858,858'b0};
assign c[2590319:2587308] = {647'b0,c_w_859,859'b0};
assign c[2593331:2590320] = {646'b0,c_w_860,860'b0};
assign c[2596343:2593332] = {645'b0,c_w_861,861'b0};
assign c[2599355:2596344] = {644'b0,c_w_862,862'b0};
assign c[2602367:2599356] = {643'b0,c_w_863,863'b0};
assign c[2605379:2602368] = {642'b0,c_w_864,864'b0};
assign c[2608391:2605380] = {641'b0,c_w_865,865'b0};
assign c[2611403:2608392] = {640'b0,c_w_866,866'b0};
assign c[2614415:2611404] = {639'b0,c_w_867,867'b0};
assign c[2617427:2614416] = {638'b0,c_w_868,868'b0};
assign c[2620439:2617428] = {637'b0,c_w_869,869'b0};
assign c[2623451:2620440] = {636'b0,c_w_870,870'b0};
assign c[2626463:2623452] = {635'b0,c_w_871,871'b0};
assign c[2629475:2626464] = {634'b0,c_w_872,872'b0};
assign c[2632487:2629476] = {633'b0,c_w_873,873'b0};
assign c[2635499:2632488] = {632'b0,c_w_874,874'b0};
assign c[2638511:2635500] = {631'b0,c_w_875,875'b0};
assign c[2641523:2638512] = {630'b0,c_w_876,876'b0};
assign c[2644535:2641524] = {629'b0,c_w_877,877'b0};
assign c[2647547:2644536] = {628'b0,c_w_878,878'b0};
assign c[2650559:2647548] = {627'b0,c_w_879,879'b0};
assign c[2653571:2650560] = {626'b0,c_w_880,880'b0};
assign c[2656583:2653572] = {625'b0,c_w_881,881'b0};
assign c[2659595:2656584] = {624'b0,c_w_882,882'b0};
assign c[2662607:2659596] = {623'b0,c_w_883,883'b0};
assign c[2665619:2662608] = {622'b0,c_w_884,884'b0};
assign c[2668631:2665620] = {621'b0,c_w_885,885'b0};
assign c[2671643:2668632] = {620'b0,c_w_886,886'b0};
assign c[2674655:2671644] = {619'b0,c_w_887,887'b0};
assign c[2677667:2674656] = {618'b0,c_w_888,888'b0};
assign c[2680679:2677668] = {617'b0,c_w_889,889'b0};
assign c[2683691:2680680] = {616'b0,c_w_890,890'b0};
assign c[2686703:2683692] = {615'b0,c_w_891,891'b0};
assign c[2689715:2686704] = {614'b0,c_w_892,892'b0};
assign c[2692727:2689716] = {613'b0,c_w_893,893'b0};
assign c[2695739:2692728] = {612'b0,c_w_894,894'b0};
assign c[2698751:2695740] = {611'b0,c_w_895,895'b0};
assign c[2701763:2698752] = {610'b0,c_w_896,896'b0};
assign c[2704775:2701764] = {609'b0,c_w_897,897'b0};
assign c[2707787:2704776] = {608'b0,c_w_898,898'b0};
assign c[2710799:2707788] = {607'b0,c_w_899,899'b0};
assign c[2713811:2710800] = {606'b0,c_w_900,900'b0};
assign c[2716823:2713812] = {605'b0,c_w_901,901'b0};
assign c[2719835:2716824] = {604'b0,c_w_902,902'b0};
assign c[2722847:2719836] = {603'b0,c_w_903,903'b0};
assign c[2725859:2722848] = {602'b0,c_w_904,904'b0};
assign c[2728871:2725860] = {601'b0,c_w_905,905'b0};
assign c[2731883:2728872] = {600'b0,c_w_906,906'b0};
assign c[2734895:2731884] = {599'b0,c_w_907,907'b0};
assign c[2737907:2734896] = {598'b0,c_w_908,908'b0};
assign c[2740919:2737908] = {597'b0,c_w_909,909'b0};
assign c[2743931:2740920] = {596'b0,c_w_910,910'b0};
assign c[2746943:2743932] = {595'b0,c_w_911,911'b0};
assign c[2749955:2746944] = {594'b0,c_w_912,912'b0};
assign c[2752967:2749956] = {593'b0,c_w_913,913'b0};
assign c[2755979:2752968] = {592'b0,c_w_914,914'b0};
assign c[2758991:2755980] = {591'b0,c_w_915,915'b0};
assign c[2762003:2758992] = {590'b0,c_w_916,916'b0};
assign c[2765015:2762004] = {589'b0,c_w_917,917'b0};
assign c[2768027:2765016] = {588'b0,c_w_918,918'b0};
assign c[2771039:2768028] = {587'b0,c_w_919,919'b0};
assign c[2774051:2771040] = {586'b0,c_w_920,920'b0};
assign c[2777063:2774052] = {585'b0,c_w_921,921'b0};
assign c[2780075:2777064] = {584'b0,c_w_922,922'b0};
assign c[2783087:2780076] = {583'b0,c_w_923,923'b0};
assign c[2786099:2783088] = {582'b0,c_w_924,924'b0};
assign c[2789111:2786100] = {581'b0,c_w_925,925'b0};
assign c[2792123:2789112] = {580'b0,c_w_926,926'b0};
assign c[2795135:2792124] = {579'b0,c_w_927,927'b0};
assign c[2798147:2795136] = {578'b0,c_w_928,928'b0};
assign c[2801159:2798148] = {577'b0,c_w_929,929'b0};
assign c[2804171:2801160] = {576'b0,c_w_930,930'b0};
assign c[2807183:2804172] = {575'b0,c_w_931,931'b0};
assign c[2810195:2807184] = {574'b0,c_w_932,932'b0};
assign c[2813207:2810196] = {573'b0,c_w_933,933'b0};
assign c[2816219:2813208] = {572'b0,c_w_934,934'b0};
assign c[2819231:2816220] = {571'b0,c_w_935,935'b0};
assign c[2822243:2819232] = {570'b0,c_w_936,936'b0};
assign c[2825255:2822244] = {569'b0,c_w_937,937'b0};
assign c[2828267:2825256] = {568'b0,c_w_938,938'b0};
assign c[2831279:2828268] = {567'b0,c_w_939,939'b0};
assign c[2834291:2831280] = {566'b0,c_w_940,940'b0};
assign c[2837303:2834292] = {565'b0,c_w_941,941'b0};
assign c[2840315:2837304] = {564'b0,c_w_942,942'b0};
assign c[2843327:2840316] = {563'b0,c_w_943,943'b0};
assign c[2846339:2843328] = {562'b0,c_w_944,944'b0};
assign c[2849351:2846340] = {561'b0,c_w_945,945'b0};
assign c[2852363:2849352] = {560'b0,c_w_946,946'b0};
assign c[2855375:2852364] = {559'b0,c_w_947,947'b0};
assign c[2858387:2855376] = {558'b0,c_w_948,948'b0};
assign c[2861399:2858388] = {557'b0,c_w_949,949'b0};
assign c[2864411:2861400] = {556'b0,c_w_950,950'b0};
assign c[2867423:2864412] = {555'b0,c_w_951,951'b0};
assign c[2870435:2867424] = {554'b0,c_w_952,952'b0};
assign c[2873447:2870436] = {553'b0,c_w_953,953'b0};
assign c[2876459:2873448] = {552'b0,c_w_954,954'b0};
assign c[2879471:2876460] = {551'b0,c_w_955,955'b0};
assign c[2882483:2879472] = {550'b0,c_w_956,956'b0};
assign c[2885495:2882484] = {549'b0,c_w_957,957'b0};
assign c[2888507:2885496] = {548'b0,c_w_958,958'b0};
assign c[2891519:2888508] = {547'b0,c_w_959,959'b0};
assign c[2894531:2891520] = {546'b0,c_w_960,960'b0};
assign c[2897543:2894532] = {545'b0,c_w_961,961'b0};
assign c[2900555:2897544] = {544'b0,c_w_962,962'b0};
assign c[2903567:2900556] = {543'b0,c_w_963,963'b0};
assign c[2906579:2903568] = {542'b0,c_w_964,964'b0};
assign c[2909591:2906580] = {541'b0,c_w_965,965'b0};
assign c[2912603:2909592] = {540'b0,c_w_966,966'b0};
assign c[2915615:2912604] = {539'b0,c_w_967,967'b0};
assign c[2918627:2915616] = {538'b0,c_w_968,968'b0};
assign c[2921639:2918628] = {537'b0,c_w_969,969'b0};
assign c[2924651:2921640] = {536'b0,c_w_970,970'b0};
assign c[2927663:2924652] = {535'b0,c_w_971,971'b0};
assign c[2930675:2927664] = {534'b0,c_w_972,972'b0};
assign c[2933687:2930676] = {533'b0,c_w_973,973'b0};
assign c[2936699:2933688] = {532'b0,c_w_974,974'b0};
assign c[2939711:2936700] = {531'b0,c_w_975,975'b0};
assign c[2942723:2939712] = {530'b0,c_w_976,976'b0};
assign c[2945735:2942724] = {529'b0,c_w_977,977'b0};
assign c[2948747:2945736] = {528'b0,c_w_978,978'b0};
assign c[2951759:2948748] = {527'b0,c_w_979,979'b0};
assign c[2954771:2951760] = {526'b0,c_w_980,980'b0};
assign c[2957783:2954772] = {525'b0,c_w_981,981'b0};
assign c[2960795:2957784] = {524'b0,c_w_982,982'b0};
assign c[2963807:2960796] = {523'b0,c_w_983,983'b0};
assign c[2966819:2963808] = {522'b0,c_w_984,984'b0};
assign c[2969831:2966820] = {521'b0,c_w_985,985'b0};
assign c[2972843:2969832] = {520'b0,c_w_986,986'b0};
assign c[2975855:2972844] = {519'b0,c_w_987,987'b0};
assign c[2978867:2975856] = {518'b0,c_w_988,988'b0};
assign c[2981879:2978868] = {517'b0,c_w_989,989'b0};
assign c[2984891:2981880] = {516'b0,c_w_990,990'b0};
assign c[2987903:2984892] = {515'b0,c_w_991,991'b0};
assign c[2990915:2987904] = {514'b0,c_w_992,992'b0};
assign c[2993927:2990916] = {513'b0,c_w_993,993'b0};
assign c[2996939:2993928] = {512'b0,c_w_994,994'b0};
assign c[2999951:2996940] = {511'b0,c_w_995,995'b0};
assign c[3002963:2999952] = {510'b0,c_w_996,996'b0};
assign c[3005975:3002964] = {509'b0,c_w_997,997'b0};
assign c[3008987:3005976] = {508'b0,c_w_998,998'b0};
assign c[3011999:3008988] = {507'b0,c_w_999,999'b0};
assign c[3015011:3012000] = {506'b0,c_w_1000,1000'b0};
assign c[3018023:3015012] = {505'b0,c_w_1001,1001'b0};
assign c[3021035:3018024] = {504'b0,c_w_1002,1002'b0};
assign c[3024047:3021036] = {503'b0,c_w_1003,1003'b0};
assign c[3027059:3024048] = {502'b0,c_w_1004,1004'b0};
assign c[3030071:3027060] = {501'b0,c_w_1005,1005'b0};
assign c[3033083:3030072] = {500'b0,c_w_1006,1006'b0};
assign c[3036095:3033084] = {499'b0,c_w_1007,1007'b0};
assign c[3039107:3036096] = {498'b0,c_w_1008,1008'b0};
assign c[3042119:3039108] = {497'b0,c_w_1009,1009'b0};
assign c[3045131:3042120] = {496'b0,c_w_1010,1010'b0};
assign c[3048143:3045132] = {495'b0,c_w_1011,1011'b0};
assign c[3051155:3048144] = {494'b0,c_w_1012,1012'b0};
assign c[3054167:3051156] = {493'b0,c_w_1013,1013'b0};
assign c[3057179:3054168] = {492'b0,c_w_1014,1014'b0};
assign c[3060191:3057180] = {491'b0,c_w_1015,1015'b0};
assign c[3063203:3060192] = {490'b0,c_w_1016,1016'b0};
assign c[3066215:3063204] = {489'b0,c_w_1017,1017'b0};
assign c[3069227:3066216] = {488'b0,c_w_1018,1018'b0};
assign c[3072239:3069228] = {487'b0,c_w_1019,1019'b0};
assign c[3075251:3072240] = {486'b0,c_w_1020,1020'b0};
assign c[3078263:3075252] = {485'b0,c_w_1021,1021'b0};
assign c[3081275:3078264] = {484'b0,c_w_1022,1022'b0};
assign c[3084287:3081276] = {483'b0,c_w_1023,1023'b0};
assign c[3087299:3084288] = {482'b0,c_w_1024,1024'b0};
assign c[3090311:3087300] = {481'b0,c_w_1025,1025'b0};
assign c[3093323:3090312] = {480'b0,c_w_1026,1026'b0};
assign c[3096335:3093324] = {479'b0,c_w_1027,1027'b0};
assign c[3099347:3096336] = {478'b0,c_w_1028,1028'b0};
assign c[3102359:3099348] = {477'b0,c_w_1029,1029'b0};
assign c[3105371:3102360] = {476'b0,c_w_1030,1030'b0};
assign c[3108383:3105372] = {475'b0,c_w_1031,1031'b0};
assign c[3111395:3108384] = {474'b0,c_w_1032,1032'b0};
assign c[3114407:3111396] = {473'b0,c_w_1033,1033'b0};
assign c[3117419:3114408] = {472'b0,c_w_1034,1034'b0};
assign c[3120431:3117420] = {471'b0,c_w_1035,1035'b0};
assign c[3123443:3120432] = {470'b0,c_w_1036,1036'b0};
assign c[3126455:3123444] = {469'b0,c_w_1037,1037'b0};
assign c[3129467:3126456] = {468'b0,c_w_1038,1038'b0};
assign c[3132479:3129468] = {467'b0,c_w_1039,1039'b0};
assign c[3135491:3132480] = {466'b0,c_w_1040,1040'b0};
assign c[3138503:3135492] = {465'b0,c_w_1041,1041'b0};
assign c[3141515:3138504] = {464'b0,c_w_1042,1042'b0};
assign c[3144527:3141516] = {463'b0,c_w_1043,1043'b0};
assign c[3147539:3144528] = {462'b0,c_w_1044,1044'b0};
assign c[3150551:3147540] = {461'b0,c_w_1045,1045'b0};
assign c[3153563:3150552] = {460'b0,c_w_1046,1046'b0};
assign c[3156575:3153564] = {459'b0,c_w_1047,1047'b0};
assign c[3159587:3156576] = {458'b0,c_w_1048,1048'b0};
assign c[3162599:3159588] = {457'b0,c_w_1049,1049'b0};
assign c[3165611:3162600] = {456'b0,c_w_1050,1050'b0};
assign c[3168623:3165612] = {455'b0,c_w_1051,1051'b0};
assign c[3171635:3168624] = {454'b0,c_w_1052,1052'b0};
assign c[3174647:3171636] = {453'b0,c_w_1053,1053'b0};
assign c[3177659:3174648] = {452'b0,c_w_1054,1054'b0};
assign c[3180671:3177660] = {451'b0,c_w_1055,1055'b0};
assign c[3183683:3180672] = {450'b0,c_w_1056,1056'b0};
assign c[3186695:3183684] = {449'b0,c_w_1057,1057'b0};
assign c[3189707:3186696] = {448'b0,c_w_1058,1058'b0};
assign c[3192719:3189708] = {447'b0,c_w_1059,1059'b0};
assign c[3195731:3192720] = {446'b0,c_w_1060,1060'b0};
assign c[3198743:3195732] = {445'b0,c_w_1061,1061'b0};
assign c[3201755:3198744] = {444'b0,c_w_1062,1062'b0};
assign c[3204767:3201756] = {443'b0,c_w_1063,1063'b0};
assign c[3207779:3204768] = {442'b0,c_w_1064,1064'b0};
assign c[3210791:3207780] = {441'b0,c_w_1065,1065'b0};
assign c[3213803:3210792] = {440'b0,c_w_1066,1066'b0};
assign c[3216815:3213804] = {439'b0,c_w_1067,1067'b0};
assign c[3219827:3216816] = {438'b0,c_w_1068,1068'b0};
assign c[3222839:3219828] = {437'b0,c_w_1069,1069'b0};
assign c[3225851:3222840] = {436'b0,c_w_1070,1070'b0};
assign c[3228863:3225852] = {435'b0,c_w_1071,1071'b0};
assign c[3231875:3228864] = {434'b0,c_w_1072,1072'b0};
assign c[3234887:3231876] = {433'b0,c_w_1073,1073'b0};
assign c[3237899:3234888] = {432'b0,c_w_1074,1074'b0};
assign c[3240911:3237900] = {431'b0,c_w_1075,1075'b0};
assign c[3243923:3240912] = {430'b0,c_w_1076,1076'b0};
assign c[3246935:3243924] = {429'b0,c_w_1077,1077'b0};
assign c[3249947:3246936] = {428'b0,c_w_1078,1078'b0};
assign c[3252959:3249948] = {427'b0,c_w_1079,1079'b0};
assign c[3255971:3252960] = {426'b0,c_w_1080,1080'b0};
assign c[3258983:3255972] = {425'b0,c_w_1081,1081'b0};
assign c[3261995:3258984] = {424'b0,c_w_1082,1082'b0};
assign c[3265007:3261996] = {423'b0,c_w_1083,1083'b0};
assign c[3268019:3265008] = {422'b0,c_w_1084,1084'b0};
assign c[3271031:3268020] = {421'b0,c_w_1085,1085'b0};
assign c[3274043:3271032] = {420'b0,c_w_1086,1086'b0};
assign c[3277055:3274044] = {419'b0,c_w_1087,1087'b0};
assign c[3280067:3277056] = {418'b0,c_w_1088,1088'b0};
assign c[3283079:3280068] = {417'b0,c_w_1089,1089'b0};
assign c[3286091:3283080] = {416'b0,c_w_1090,1090'b0};
assign c[3289103:3286092] = {415'b0,c_w_1091,1091'b0};
assign c[3292115:3289104] = {414'b0,c_w_1092,1092'b0};
assign c[3295127:3292116] = {413'b0,c_w_1093,1093'b0};
assign c[3298139:3295128] = {412'b0,c_w_1094,1094'b0};
assign c[3301151:3298140] = {411'b0,c_w_1095,1095'b0};
assign c[3304163:3301152] = {410'b0,c_w_1096,1096'b0};
assign c[3307175:3304164] = {409'b0,c_w_1097,1097'b0};
assign c[3310187:3307176] = {408'b0,c_w_1098,1098'b0};
assign c[3313199:3310188] = {407'b0,c_w_1099,1099'b0};
assign c[3316211:3313200] = {406'b0,c_w_1100,1100'b0};
assign c[3319223:3316212] = {405'b0,c_w_1101,1101'b0};
assign c[3322235:3319224] = {404'b0,c_w_1102,1102'b0};
assign c[3325247:3322236] = {403'b0,c_w_1103,1103'b0};
assign c[3328259:3325248] = {402'b0,c_w_1104,1104'b0};
assign c[3331271:3328260] = {401'b0,c_w_1105,1105'b0};
assign c[3334283:3331272] = {400'b0,c_w_1106,1106'b0};
assign c[3337295:3334284] = {399'b0,c_w_1107,1107'b0};
assign c[3340307:3337296] = {398'b0,c_w_1108,1108'b0};
assign c[3343319:3340308] = {397'b0,c_w_1109,1109'b0};
assign c[3346331:3343320] = {396'b0,c_w_1110,1110'b0};
assign c[3349343:3346332] = {395'b0,c_w_1111,1111'b0};
assign c[3352355:3349344] = {394'b0,c_w_1112,1112'b0};
assign c[3355367:3352356] = {393'b0,c_w_1113,1113'b0};
assign c[3358379:3355368] = {392'b0,c_w_1114,1114'b0};
assign c[3361391:3358380] = {391'b0,c_w_1115,1115'b0};
assign c[3364403:3361392] = {390'b0,c_w_1116,1116'b0};
assign c[3367415:3364404] = {389'b0,c_w_1117,1117'b0};
assign c[3370427:3367416] = {388'b0,c_w_1118,1118'b0};
assign c[3373439:3370428] = {387'b0,c_w_1119,1119'b0};
assign c[3376451:3373440] = {386'b0,c_w_1120,1120'b0};
assign c[3379463:3376452] = {385'b0,c_w_1121,1121'b0};
assign c[3382475:3379464] = {384'b0,c_w_1122,1122'b0};
assign c[3385487:3382476] = {383'b0,c_w_1123,1123'b0};
assign c[3388499:3385488] = {382'b0,c_w_1124,1124'b0};
assign c[3391511:3388500] = {381'b0,c_w_1125,1125'b0};
assign c[3394523:3391512] = {380'b0,c_w_1126,1126'b0};
assign c[3397535:3394524] = {379'b0,c_w_1127,1127'b0};
assign c[3400547:3397536] = {378'b0,c_w_1128,1128'b0};
assign c[3403559:3400548] = {377'b0,c_w_1129,1129'b0};
assign c[3406571:3403560] = {376'b0,c_w_1130,1130'b0};
assign c[3409583:3406572] = {375'b0,c_w_1131,1131'b0};
assign c[3412595:3409584] = {374'b0,c_w_1132,1132'b0};
assign c[3415607:3412596] = {373'b0,c_w_1133,1133'b0};
assign c[3418619:3415608] = {372'b0,c_w_1134,1134'b0};
assign c[3421631:3418620] = {371'b0,c_w_1135,1135'b0};
assign c[3424643:3421632] = {370'b0,c_w_1136,1136'b0};
assign c[3427655:3424644] = {369'b0,c_w_1137,1137'b0};
assign c[3430667:3427656] = {368'b0,c_w_1138,1138'b0};
assign c[3433679:3430668] = {367'b0,c_w_1139,1139'b0};
assign c[3436691:3433680] = {366'b0,c_w_1140,1140'b0};
assign c[3439703:3436692] = {365'b0,c_w_1141,1141'b0};
assign c[3442715:3439704] = {364'b0,c_w_1142,1142'b0};
assign c[3445727:3442716] = {363'b0,c_w_1143,1143'b0};
assign c[3448739:3445728] = {362'b0,c_w_1144,1144'b0};
assign c[3451751:3448740] = {361'b0,c_w_1145,1145'b0};
assign c[3454763:3451752] = {360'b0,c_w_1146,1146'b0};
assign c[3457775:3454764] = {359'b0,c_w_1147,1147'b0};
assign c[3460787:3457776] = {358'b0,c_w_1148,1148'b0};
assign c[3463799:3460788] = {357'b0,c_w_1149,1149'b0};
assign c[3466811:3463800] = {356'b0,c_w_1150,1150'b0};
assign c[3469823:3466812] = {355'b0,c_w_1151,1151'b0};
assign c[3472835:3469824] = {354'b0,c_w_1152,1152'b0};
assign c[3475847:3472836] = {353'b0,c_w_1153,1153'b0};
assign c[3478859:3475848] = {352'b0,c_w_1154,1154'b0};
assign c[3481871:3478860] = {351'b0,c_w_1155,1155'b0};
assign c[3484883:3481872] = {350'b0,c_w_1156,1156'b0};
assign c[3487895:3484884] = {349'b0,c_w_1157,1157'b0};
assign c[3490907:3487896] = {348'b0,c_w_1158,1158'b0};
assign c[3493919:3490908] = {347'b0,c_w_1159,1159'b0};
assign c[3496931:3493920] = {346'b0,c_w_1160,1160'b0};
assign c[3499943:3496932] = {345'b0,c_w_1161,1161'b0};
assign c[3502955:3499944] = {344'b0,c_w_1162,1162'b0};
assign c[3505967:3502956] = {343'b0,c_w_1163,1163'b0};
assign c[3508979:3505968] = {342'b0,c_w_1164,1164'b0};
assign c[3511991:3508980] = {341'b0,c_w_1165,1165'b0};
assign c[3515003:3511992] = {340'b0,c_w_1166,1166'b0};
assign c[3518015:3515004] = {339'b0,c_w_1167,1167'b0};
assign c[3521027:3518016] = {338'b0,c_w_1168,1168'b0};
assign c[3524039:3521028] = {337'b0,c_w_1169,1169'b0};
assign c[3527051:3524040] = {336'b0,c_w_1170,1170'b0};
assign c[3530063:3527052] = {335'b0,c_w_1171,1171'b0};
assign c[3533075:3530064] = {334'b0,c_w_1172,1172'b0};
assign c[3536087:3533076] = {333'b0,c_w_1173,1173'b0};
assign c[3539099:3536088] = {332'b0,c_w_1174,1174'b0};
assign c[3542111:3539100] = {331'b0,c_w_1175,1175'b0};
assign c[3545123:3542112] = {330'b0,c_w_1176,1176'b0};
assign c[3548135:3545124] = {329'b0,c_w_1177,1177'b0};
assign c[3551147:3548136] = {328'b0,c_w_1178,1178'b0};
assign c[3554159:3551148] = {327'b0,c_w_1179,1179'b0};
assign c[3557171:3554160] = {326'b0,c_w_1180,1180'b0};
assign c[3560183:3557172] = {325'b0,c_w_1181,1181'b0};
assign c[3563195:3560184] = {324'b0,c_w_1182,1182'b0};
assign c[3566207:3563196] = {323'b0,c_w_1183,1183'b0};
assign c[3569219:3566208] = {322'b0,c_w_1184,1184'b0};
assign c[3572231:3569220] = {321'b0,c_w_1185,1185'b0};
assign c[3575243:3572232] = {320'b0,c_w_1186,1186'b0};
assign c[3578255:3575244] = {319'b0,c_w_1187,1187'b0};
assign c[3581267:3578256] = {318'b0,c_w_1188,1188'b0};
assign c[3584279:3581268] = {317'b0,c_w_1189,1189'b0};
assign c[3587291:3584280] = {316'b0,c_w_1190,1190'b0};
assign c[3590303:3587292] = {315'b0,c_w_1191,1191'b0};
assign c[3593315:3590304] = {314'b0,c_w_1192,1192'b0};
assign c[3596327:3593316] = {313'b0,c_w_1193,1193'b0};
assign c[3599339:3596328] = {312'b0,c_w_1194,1194'b0};
assign c[3602351:3599340] = {311'b0,c_w_1195,1195'b0};
assign c[3605363:3602352] = {310'b0,c_w_1196,1196'b0};
assign c[3608375:3605364] = {309'b0,c_w_1197,1197'b0};
assign c[3611387:3608376] = {308'b0,c_w_1198,1198'b0};
assign c[3614399:3611388] = {307'b0,c_w_1199,1199'b0};
assign c[3617411:3614400] = {306'b0,c_w_1200,1200'b0};
assign c[3620423:3617412] = {305'b0,c_w_1201,1201'b0};
assign c[3623435:3620424] = {304'b0,c_w_1202,1202'b0};
assign c[3626447:3623436] = {303'b0,c_w_1203,1203'b0};
assign c[3629459:3626448] = {302'b0,c_w_1204,1204'b0};
assign c[3632471:3629460] = {301'b0,c_w_1205,1205'b0};
assign c[3635483:3632472] = {300'b0,c_w_1206,1206'b0};
assign c[3638495:3635484] = {299'b0,c_w_1207,1207'b0};
assign c[3641507:3638496] = {298'b0,c_w_1208,1208'b0};
assign c[3644519:3641508] = {297'b0,c_w_1209,1209'b0};
assign c[3647531:3644520] = {296'b0,c_w_1210,1210'b0};
assign c[3650543:3647532] = {295'b0,c_w_1211,1211'b0};
assign c[3653555:3650544] = {294'b0,c_w_1212,1212'b0};
assign c[3656567:3653556] = {293'b0,c_w_1213,1213'b0};
assign c[3659579:3656568] = {292'b0,c_w_1214,1214'b0};
assign c[3662591:3659580] = {291'b0,c_w_1215,1215'b0};
assign c[3665603:3662592] = {290'b0,c_w_1216,1216'b0};
assign c[3668615:3665604] = {289'b0,c_w_1217,1217'b0};
assign c[3671627:3668616] = {288'b0,c_w_1218,1218'b0};
assign c[3674639:3671628] = {287'b0,c_w_1219,1219'b0};
assign c[3677651:3674640] = {286'b0,c_w_1220,1220'b0};
assign c[3680663:3677652] = {285'b0,c_w_1221,1221'b0};
assign c[3683675:3680664] = {284'b0,c_w_1222,1222'b0};
assign c[3686687:3683676] = {283'b0,c_w_1223,1223'b0};
assign c[3689699:3686688] = {282'b0,c_w_1224,1224'b0};
assign c[3692711:3689700] = {281'b0,c_w_1225,1225'b0};
assign c[3695723:3692712] = {280'b0,c_w_1226,1226'b0};
assign c[3698735:3695724] = {279'b0,c_w_1227,1227'b0};
assign c[3701747:3698736] = {278'b0,c_w_1228,1228'b0};
assign c[3704759:3701748] = {277'b0,c_w_1229,1229'b0};
assign c[3707771:3704760] = {276'b0,c_w_1230,1230'b0};
assign c[3710783:3707772] = {275'b0,c_w_1231,1231'b0};
assign c[3713795:3710784] = {274'b0,c_w_1232,1232'b0};
assign c[3716807:3713796] = {273'b0,c_w_1233,1233'b0};
assign c[3719819:3716808] = {272'b0,c_w_1234,1234'b0};
assign c[3722831:3719820] = {271'b0,c_w_1235,1235'b0};
assign c[3725843:3722832] = {270'b0,c_w_1236,1236'b0};
assign c[3728855:3725844] = {269'b0,c_w_1237,1237'b0};
assign c[3731867:3728856] = {268'b0,c_w_1238,1238'b0};
assign c[3734879:3731868] = {267'b0,c_w_1239,1239'b0};
assign c[3737891:3734880] = {266'b0,c_w_1240,1240'b0};
assign c[3740903:3737892] = {265'b0,c_w_1241,1241'b0};
assign c[3743915:3740904] = {264'b0,c_w_1242,1242'b0};
assign c[3746927:3743916] = {263'b0,c_w_1243,1243'b0};
assign c[3749939:3746928] = {262'b0,c_w_1244,1244'b0};
assign c[3752951:3749940] = {261'b0,c_w_1245,1245'b0};
assign c[3755963:3752952] = {260'b0,c_w_1246,1246'b0};
assign c[3758975:3755964] = {259'b0,c_w_1247,1247'b0};
assign c[3761987:3758976] = {258'b0,c_w_1248,1248'b0};
assign c[3764999:3761988] = {257'b0,c_w_1249,1249'b0};
assign c[3768011:3765000] = {256'b0,c_w_1250,1250'b0};
assign c[3771023:3768012] = {255'b0,c_w_1251,1251'b0};
assign c[3774035:3771024] = {254'b0,c_w_1252,1252'b0};
assign c[3777047:3774036] = {253'b0,c_w_1253,1253'b0};
assign c[3780059:3777048] = {252'b0,c_w_1254,1254'b0};
assign c[3783071:3780060] = {251'b0,c_w_1255,1255'b0};
assign c[3786083:3783072] = {250'b0,c_w_1256,1256'b0};
assign c[3789095:3786084] = {249'b0,c_w_1257,1257'b0};
assign c[3792107:3789096] = {248'b0,c_w_1258,1258'b0};
assign c[3795119:3792108] = {247'b0,c_w_1259,1259'b0};
assign c[3798131:3795120] = {246'b0,c_w_1260,1260'b0};
assign c[3801143:3798132] = {245'b0,c_w_1261,1261'b0};
assign c[3804155:3801144] = {244'b0,c_w_1262,1262'b0};
assign c[3807167:3804156] = {243'b0,c_w_1263,1263'b0};
assign c[3810179:3807168] = {242'b0,c_w_1264,1264'b0};
assign c[3813191:3810180] = {241'b0,c_w_1265,1265'b0};
assign c[3816203:3813192] = {240'b0,c_w_1266,1266'b0};
assign c[3819215:3816204] = {239'b0,c_w_1267,1267'b0};
assign c[3822227:3819216] = {238'b0,c_w_1268,1268'b0};
assign c[3825239:3822228] = {237'b0,c_w_1269,1269'b0};
assign c[3828251:3825240] = {236'b0,c_w_1270,1270'b0};
assign c[3831263:3828252] = {235'b0,c_w_1271,1271'b0};
assign c[3834275:3831264] = {234'b0,c_w_1272,1272'b0};
assign c[3837287:3834276] = {233'b0,c_w_1273,1273'b0};
assign c[3840299:3837288] = {232'b0,c_w_1274,1274'b0};
assign c[3843311:3840300] = {231'b0,c_w_1275,1275'b0};
assign c[3846323:3843312] = {230'b0,c_w_1276,1276'b0};
assign c[3849335:3846324] = {229'b0,c_w_1277,1277'b0};
assign c[3852347:3849336] = {228'b0,c_w_1278,1278'b0};
assign c[3855359:3852348] = {227'b0,c_w_1279,1279'b0};
assign c[3858371:3855360] = {226'b0,c_w_1280,1280'b0};
assign c[3861383:3858372] = {225'b0,c_w_1281,1281'b0};
assign c[3864395:3861384] = {224'b0,c_w_1282,1282'b0};
assign c[3867407:3864396] = {223'b0,c_w_1283,1283'b0};
assign c[3870419:3867408] = {222'b0,c_w_1284,1284'b0};
assign c[3873431:3870420] = {221'b0,c_w_1285,1285'b0};
assign c[3876443:3873432] = {220'b0,c_w_1286,1286'b0};
assign c[3879455:3876444] = {219'b0,c_w_1287,1287'b0};
assign c[3882467:3879456] = {218'b0,c_w_1288,1288'b0};
assign c[3885479:3882468] = {217'b0,c_w_1289,1289'b0};
assign c[3888491:3885480] = {216'b0,c_w_1290,1290'b0};
assign c[3891503:3888492] = {215'b0,c_w_1291,1291'b0};
assign c[3894515:3891504] = {214'b0,c_w_1292,1292'b0};
assign c[3897527:3894516] = {213'b0,c_w_1293,1293'b0};
assign c[3900539:3897528] = {212'b0,c_w_1294,1294'b0};
assign c[3903551:3900540] = {211'b0,c_w_1295,1295'b0};
assign c[3906563:3903552] = {210'b0,c_w_1296,1296'b0};
assign c[3909575:3906564] = {209'b0,c_w_1297,1297'b0};
assign c[3912587:3909576] = {208'b0,c_w_1298,1298'b0};
assign c[3915599:3912588] = {207'b0,c_w_1299,1299'b0};
assign c[3918611:3915600] = {206'b0,c_w_1300,1300'b0};
assign c[3921623:3918612] = {205'b0,c_w_1301,1301'b0};
assign c[3924635:3921624] = {204'b0,c_w_1302,1302'b0};
assign c[3927647:3924636] = {203'b0,c_w_1303,1303'b0};
assign c[3930659:3927648] = {202'b0,c_w_1304,1304'b0};
assign c[3933671:3930660] = {201'b0,c_w_1305,1305'b0};
assign c[3936683:3933672] = {200'b0,c_w_1306,1306'b0};
assign c[3939695:3936684] = {199'b0,c_w_1307,1307'b0};
assign c[3942707:3939696] = {198'b0,c_w_1308,1308'b0};
assign c[3945719:3942708] = {197'b0,c_w_1309,1309'b0};
assign c[3948731:3945720] = {196'b0,c_w_1310,1310'b0};
assign c[3951743:3948732] = {195'b0,c_w_1311,1311'b0};
assign c[3954755:3951744] = {194'b0,c_w_1312,1312'b0};
assign c[3957767:3954756] = {193'b0,c_w_1313,1313'b0};
assign c[3960779:3957768] = {192'b0,c_w_1314,1314'b0};
assign c[3963791:3960780] = {191'b0,c_w_1315,1315'b0};
assign c[3966803:3963792] = {190'b0,c_w_1316,1316'b0};
assign c[3969815:3966804] = {189'b0,c_w_1317,1317'b0};
assign c[3972827:3969816] = {188'b0,c_w_1318,1318'b0};
assign c[3975839:3972828] = {187'b0,c_w_1319,1319'b0};
assign c[3978851:3975840] = {186'b0,c_w_1320,1320'b0};
assign c[3981863:3978852] = {185'b0,c_w_1321,1321'b0};
assign c[3984875:3981864] = {184'b0,c_w_1322,1322'b0};
assign c[3987887:3984876] = {183'b0,c_w_1323,1323'b0};
assign c[3990899:3987888] = {182'b0,c_w_1324,1324'b0};
assign c[3993911:3990900] = {181'b0,c_w_1325,1325'b0};
assign c[3996923:3993912] = {180'b0,c_w_1326,1326'b0};
assign c[3999935:3996924] = {179'b0,c_w_1327,1327'b0};
assign c[4002947:3999936] = {178'b0,c_w_1328,1328'b0};
assign c[4005959:4002948] = {177'b0,c_w_1329,1329'b0};
assign c[4008971:4005960] = {176'b0,c_w_1330,1330'b0};
assign c[4011983:4008972] = {175'b0,c_w_1331,1331'b0};
assign c[4014995:4011984] = {174'b0,c_w_1332,1332'b0};
assign c[4018007:4014996] = {173'b0,c_w_1333,1333'b0};
assign c[4021019:4018008] = {172'b0,c_w_1334,1334'b0};
assign c[4024031:4021020] = {171'b0,c_w_1335,1335'b0};
assign c[4027043:4024032] = {170'b0,c_w_1336,1336'b0};
assign c[4030055:4027044] = {169'b0,c_w_1337,1337'b0};
assign c[4033067:4030056] = {168'b0,c_w_1338,1338'b0};
assign c[4036079:4033068] = {167'b0,c_w_1339,1339'b0};
assign c[4039091:4036080] = {166'b0,c_w_1340,1340'b0};
assign c[4042103:4039092] = {165'b0,c_w_1341,1341'b0};
assign c[4045115:4042104] = {164'b0,c_w_1342,1342'b0};
assign c[4048127:4045116] = {163'b0,c_w_1343,1343'b0};
assign c[4051139:4048128] = {162'b0,c_w_1344,1344'b0};
assign c[4054151:4051140] = {161'b0,c_w_1345,1345'b0};
assign c[4057163:4054152] = {160'b0,c_w_1346,1346'b0};
assign c[4060175:4057164] = {159'b0,c_w_1347,1347'b0};
assign c[4063187:4060176] = {158'b0,c_w_1348,1348'b0};
assign c[4066199:4063188] = {157'b0,c_w_1349,1349'b0};
assign c[4069211:4066200] = {156'b0,c_w_1350,1350'b0};
assign c[4072223:4069212] = {155'b0,c_w_1351,1351'b0};
assign c[4075235:4072224] = {154'b0,c_w_1352,1352'b0};
assign c[4078247:4075236] = {153'b0,c_w_1353,1353'b0};
assign c[4081259:4078248] = {152'b0,c_w_1354,1354'b0};
assign c[4084271:4081260] = {151'b0,c_w_1355,1355'b0};
assign c[4087283:4084272] = {150'b0,c_w_1356,1356'b0};
assign c[4090295:4087284] = {149'b0,c_w_1357,1357'b0};
assign c[4093307:4090296] = {148'b0,c_w_1358,1358'b0};
assign c[4096319:4093308] = {147'b0,c_w_1359,1359'b0};
assign c[4099331:4096320] = {146'b0,c_w_1360,1360'b0};
assign c[4102343:4099332] = {145'b0,c_w_1361,1361'b0};
assign c[4105355:4102344] = {144'b0,c_w_1362,1362'b0};
assign c[4108367:4105356] = {143'b0,c_w_1363,1363'b0};
assign c[4111379:4108368] = {142'b0,c_w_1364,1364'b0};
assign c[4114391:4111380] = {141'b0,c_w_1365,1365'b0};
assign c[4117403:4114392] = {140'b0,c_w_1366,1366'b0};
assign c[4120415:4117404] = {139'b0,c_w_1367,1367'b0};
assign c[4123427:4120416] = {138'b0,c_w_1368,1368'b0};
assign c[4126439:4123428] = {137'b0,c_w_1369,1369'b0};
assign c[4129451:4126440] = {136'b0,c_w_1370,1370'b0};
assign c[4132463:4129452] = {135'b0,c_w_1371,1371'b0};
assign c[4135475:4132464] = {134'b0,c_w_1372,1372'b0};
assign c[4138487:4135476] = {133'b0,c_w_1373,1373'b0};
assign c[4141499:4138488] = {132'b0,c_w_1374,1374'b0};
assign c[4144511:4141500] = {131'b0,c_w_1375,1375'b0};
assign c[4147523:4144512] = {130'b0,c_w_1376,1376'b0};
assign c[4150535:4147524] = {129'b0,c_w_1377,1377'b0};
assign c[4153547:4150536] = {128'b0,c_w_1378,1378'b0};
assign c[4156559:4153548] = {127'b0,c_w_1379,1379'b0};
assign c[4159571:4156560] = {126'b0,c_w_1380,1380'b0};
assign c[4162583:4159572] = {125'b0,c_w_1381,1381'b0};
assign c[4165595:4162584] = {124'b0,c_w_1382,1382'b0};
assign c[4168607:4165596] = {123'b0,c_w_1383,1383'b0};
assign c[4171619:4168608] = {122'b0,c_w_1384,1384'b0};
assign c[4174631:4171620] = {121'b0,c_w_1385,1385'b0};
assign c[4177643:4174632] = {120'b0,c_w_1386,1386'b0};
assign c[4180655:4177644] = {119'b0,c_w_1387,1387'b0};
assign c[4183667:4180656] = {118'b0,c_w_1388,1388'b0};
assign c[4186679:4183668] = {117'b0,c_w_1389,1389'b0};
assign c[4189691:4186680] = {116'b0,c_w_1390,1390'b0};
assign c[4192703:4189692] = {115'b0,c_w_1391,1391'b0};
assign c[4195715:4192704] = {114'b0,c_w_1392,1392'b0};
assign c[4198727:4195716] = {113'b0,c_w_1393,1393'b0};
assign c[4201739:4198728] = {112'b0,c_w_1394,1394'b0};
assign c[4204751:4201740] = {111'b0,c_w_1395,1395'b0};
assign c[4207763:4204752] = {110'b0,c_w_1396,1396'b0};
assign c[4210775:4207764] = {109'b0,c_w_1397,1397'b0};
assign c[4213787:4210776] = {108'b0,c_w_1398,1398'b0};
assign c[4216799:4213788] = {107'b0,c_w_1399,1399'b0};
assign c[4219811:4216800] = {106'b0,c_w_1400,1400'b0};
assign c[4222823:4219812] = {105'b0,c_w_1401,1401'b0};
assign c[4225835:4222824] = {104'b0,c_w_1402,1402'b0};
assign c[4228847:4225836] = {103'b0,c_w_1403,1403'b0};
assign c[4231859:4228848] = {102'b0,c_w_1404,1404'b0};
assign c[4234871:4231860] = {101'b0,c_w_1405,1405'b0};
assign c[4237883:4234872] = {100'b0,c_w_1406,1406'b0};
assign c[4240895:4237884] = {99'b0,c_w_1407,1407'b0};
assign c[4243907:4240896] = {98'b0,c_w_1408,1408'b0};
assign c[4246919:4243908] = {97'b0,c_w_1409,1409'b0};
assign c[4249931:4246920] = {96'b0,c_w_1410,1410'b0};
assign c[4252943:4249932] = {95'b0,c_w_1411,1411'b0};
assign c[4255955:4252944] = {94'b0,c_w_1412,1412'b0};
assign c[4258967:4255956] = {93'b0,c_w_1413,1413'b0};
assign c[4261979:4258968] = {92'b0,c_w_1414,1414'b0};
assign c[4264991:4261980] = {91'b0,c_w_1415,1415'b0};
assign c[4268003:4264992] = {90'b0,c_w_1416,1416'b0};
assign c[4271015:4268004] = {89'b0,c_w_1417,1417'b0};
assign c[4274027:4271016] = {88'b0,c_w_1418,1418'b0};
assign c[4277039:4274028] = {87'b0,c_w_1419,1419'b0};
assign c[4280051:4277040] = {86'b0,c_w_1420,1420'b0};
assign c[4283063:4280052] = {85'b0,c_w_1421,1421'b0};
assign c[4286075:4283064] = {84'b0,c_w_1422,1422'b0};
assign c[4289087:4286076] = {83'b0,c_w_1423,1423'b0};
assign c[4292099:4289088] = {82'b0,c_w_1424,1424'b0};
assign c[4295111:4292100] = {81'b0,c_w_1425,1425'b0};
assign c[4298123:4295112] = {80'b0,c_w_1426,1426'b0};
assign c[4301135:4298124] = {79'b0,c_w_1427,1427'b0};
assign c[4304147:4301136] = {78'b0,c_w_1428,1428'b0};
assign c[4307159:4304148] = {77'b0,c_w_1429,1429'b0};
assign c[4310171:4307160] = {76'b0,c_w_1430,1430'b0};
assign c[4313183:4310172] = {75'b0,c_w_1431,1431'b0};
assign c[4316195:4313184] = {74'b0,c_w_1432,1432'b0};
assign c[4319207:4316196] = {73'b0,c_w_1433,1433'b0};
assign c[4322219:4319208] = {72'b0,c_w_1434,1434'b0};
assign c[4325231:4322220] = {71'b0,c_w_1435,1435'b0};
assign c[4328243:4325232] = {70'b0,c_w_1436,1436'b0};
assign c[4331255:4328244] = {69'b0,c_w_1437,1437'b0};
assign c[4334267:4331256] = {68'b0,c_w_1438,1438'b0};
assign c[4337279:4334268] = {67'b0,c_w_1439,1439'b0};
assign c[4340291:4337280] = {66'b0,c_w_1440,1440'b0};
assign c[4343303:4340292] = {65'b0,c_w_1441,1441'b0};
assign c[4346315:4343304] = {64'b0,c_w_1442,1442'b0};
assign c[4349327:4346316] = {63'b0,c_w_1443,1443'b0};
assign c[4352339:4349328] = {62'b0,c_w_1444,1444'b0};
assign c[4355351:4352340] = {61'b0,c_w_1445,1445'b0};
assign c[4358363:4355352] = {60'b0,c_w_1446,1446'b0};
assign c[4361375:4358364] = {59'b0,c_w_1447,1447'b0};
assign c[4364387:4361376] = {58'b0,c_w_1448,1448'b0};
assign c[4367399:4364388] = {57'b0,c_w_1449,1449'b0};
assign c[4370411:4367400] = {56'b0,c_w_1450,1450'b0};
assign c[4373423:4370412] = {55'b0,c_w_1451,1451'b0};
assign c[4376435:4373424] = {54'b0,c_w_1452,1452'b0};
assign c[4379447:4376436] = {53'b0,c_w_1453,1453'b0};
assign c[4382459:4379448] = {52'b0,c_w_1454,1454'b0};
assign c[4385471:4382460] = {51'b0,c_w_1455,1455'b0};
assign c[4388483:4385472] = {50'b0,c_w_1456,1456'b0};
assign c[4391495:4388484] = {49'b0,c_w_1457,1457'b0};
assign c[4394507:4391496] = {48'b0,c_w_1458,1458'b0};
assign c[4397519:4394508] = {47'b0,c_w_1459,1459'b0};
assign c[4400531:4397520] = {46'b0,c_w_1460,1460'b0};
assign c[4403543:4400532] = {45'b0,c_w_1461,1461'b0};
assign c[4406555:4403544] = {44'b0,c_w_1462,1462'b0};
assign c[4409567:4406556] = {43'b0,c_w_1463,1463'b0};
assign c[4412579:4409568] = {42'b0,c_w_1464,1464'b0};
assign c[4415591:4412580] = {41'b0,c_w_1465,1465'b0};
assign c[4418603:4415592] = {40'b0,c_w_1466,1466'b0};
assign c[4421615:4418604] = {39'b0,c_w_1467,1467'b0};
assign c[4424627:4421616] = {38'b0,c_w_1468,1468'b0};
assign c[4427639:4424628] = {37'b0,c_w_1469,1469'b0};
assign c[4430651:4427640] = {36'b0,c_w_1470,1470'b0};
assign c[4433663:4430652] = {35'b0,c_w_1471,1471'b0};
assign c[4436675:4433664] = {34'b0,c_w_1472,1472'b0};
assign c[4439687:4436676] = {33'b0,c_w_1473,1473'b0};
assign c[4442699:4439688] = {32'b0,c_w_1474,1474'b0};
assign c[4445711:4442700] = {31'b0,c_w_1475,1475'b0};
assign c[4448723:4445712] = {30'b0,c_w_1476,1476'b0};
assign c[4451735:4448724] = {29'b0,c_w_1477,1477'b0};
assign c[4454747:4451736] = {28'b0,c_w_1478,1478'b0};
assign c[4457759:4454748] = {27'b0,c_w_1479,1479'b0};
assign c[4460771:4457760] = {26'b0,c_w_1480,1480'b0};
assign c[4463783:4460772] = {25'b0,c_w_1481,1481'b0};
assign c[4466795:4463784] = {24'b0,c_w_1482,1482'b0};
assign c[4469807:4466796] = {23'b0,c_w_1483,1483'b0};
assign c[4472819:4469808] = {22'b0,c_w_1484,1484'b0};
assign c[4475831:4472820] = {21'b0,c_w_1485,1485'b0};
assign c[4478843:4475832] = {20'b0,c_w_1486,1486'b0};
assign c[4481855:4478844] = {19'b0,c_w_1487,1487'b0};
assign c[4484867:4481856] = {18'b0,c_w_1488,1488'b0};
assign c[4487879:4484868] = {17'b0,c_w_1489,1489'b0};
assign c[4490891:4487880] = {16'b0,c_w_1490,1490'b0};
assign c[4493903:4490892] = {15'b0,c_w_1491,1491'b0};
assign c[4496915:4493904] = {14'b0,c_w_1492,1492'b0};
assign c[4499927:4496916] = {13'b0,c_w_1493,1493'b0};
assign c[4502939:4499928] = {12'b0,c_w_1494,1494'b0};
assign c[4505951:4502940] = {11'b0,c_w_1495,1495'b0};
assign c[4508963:4505952] = {10'b0,c_w_1496,1496'b0};
assign c[4511975:4508964] = {9'b0,c_w_1497,1497'b0};
assign c[4514987:4511976] = {8'b0,c_w_1498,1498'b0};
assign c[4517999:4514988] = {7'b0,c_w_1499,1499'b0};
assign c[4521011:4518000] = {6'b0,c_w_1500,1500'b0};
assign c[4524023:4521012] = {5'b0,c_w_1501,1501'b0};
assign c[4527035:4524024] = {4'b0,c_w_1502,1502'b0};
assign c[4530047:4527036] = {3'b0,c_w_1503,1503'b0};
assign c[4533059:4530048] = {2'b0,c_w_1504,1504'b0};
assign c[4536071:4533060] = {1'b0,c_w_1505,1505'b0};
    
endmodule
    