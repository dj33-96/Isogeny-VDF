
module csa_186 (
    input [185:0] x,y,z,
    output[185:0] c,s 
);

wire dummy;

assign c[0] = 1'b0;
    
assign {c[1],s[0]} = (x[0]+y[0]+z[0]);
assign {c[2],s[1]} = (x[1]+y[1]+z[1]);
assign {c[3],s[2]} = (x[2]+y[2]+z[2]);
assign {c[4],s[3]} = (x[3]+y[3]+z[3]);
assign {c[5],s[4]} = (x[4]+y[4]+z[4]);
assign {c[6],s[5]} = (x[5]+y[5]+z[5]);
assign {c[7],s[6]} = (x[6]+y[6]+z[6]);
assign {c[8],s[7]} = (x[7]+y[7]+z[7]);
assign {c[9],s[8]} = (x[8]+y[8]+z[8]);
assign {c[10],s[9]} = (x[9]+y[9]+z[9]);
assign {c[11],s[10]} = (x[10]+y[10]+z[10]);
assign {c[12],s[11]} = (x[11]+y[11]+z[11]);
assign {c[13],s[12]} = (x[12]+y[12]+z[12]);
assign {c[14],s[13]} = (x[13]+y[13]+z[13]);
assign {c[15],s[14]} = (x[14]+y[14]+z[14]);
assign {c[16],s[15]} = (x[15]+y[15]+z[15]);
assign {c[17],s[16]} = (x[16]+y[16]+z[16]);
assign {c[18],s[17]} = (x[17]+y[17]+z[17]);
assign {c[19],s[18]} = (x[18]+y[18]+z[18]);
assign {c[20],s[19]} = (x[19]+y[19]+z[19]);
assign {c[21],s[20]} = (x[20]+y[20]+z[20]);
assign {c[22],s[21]} = (x[21]+y[21]+z[21]);
assign {c[23],s[22]} = (x[22]+y[22]+z[22]);
assign {c[24],s[23]} = (x[23]+y[23]+z[23]);
assign {c[25],s[24]} = (x[24]+y[24]+z[24]);
assign {c[26],s[25]} = (x[25]+y[25]+z[25]);
assign {c[27],s[26]} = (x[26]+y[26]+z[26]);
assign {c[28],s[27]} = (x[27]+y[27]+z[27]);
assign {c[29],s[28]} = (x[28]+y[28]+z[28]);
assign {c[30],s[29]} = (x[29]+y[29]+z[29]);
assign {c[31],s[30]} = (x[30]+y[30]+z[30]);
assign {c[32],s[31]} = (x[31]+y[31]+z[31]);
assign {c[33],s[32]} = (x[32]+y[32]+z[32]);
assign {c[34],s[33]} = (x[33]+y[33]+z[33]);
assign {c[35],s[34]} = (x[34]+y[34]+z[34]);
assign {c[36],s[35]} = (x[35]+y[35]+z[35]);
assign {c[37],s[36]} = (x[36]+y[36]+z[36]);
assign {c[38],s[37]} = (x[37]+y[37]+z[37]);
assign {c[39],s[38]} = (x[38]+y[38]+z[38]);
assign {c[40],s[39]} = (x[39]+y[39]+z[39]);
assign {c[41],s[40]} = (x[40]+y[40]+z[40]);
assign {c[42],s[41]} = (x[41]+y[41]+z[41]);
assign {c[43],s[42]} = (x[42]+y[42]+z[42]);
assign {c[44],s[43]} = (x[43]+y[43]+z[43]);
assign {c[45],s[44]} = (x[44]+y[44]+z[44]);
assign {c[46],s[45]} = (x[45]+y[45]+z[45]);
assign {c[47],s[46]} = (x[46]+y[46]+z[46]);
assign {c[48],s[47]} = (x[47]+y[47]+z[47]);
assign {c[49],s[48]} = (x[48]+y[48]+z[48]);
assign {c[50],s[49]} = (x[49]+y[49]+z[49]);
assign {c[51],s[50]} = (x[50]+y[50]+z[50]);
assign {c[52],s[51]} = (x[51]+y[51]+z[51]);
assign {c[53],s[52]} = (x[52]+y[52]+z[52]);
assign {c[54],s[53]} = (x[53]+y[53]+z[53]);
assign {c[55],s[54]} = (x[54]+y[54]+z[54]);
assign {c[56],s[55]} = (x[55]+y[55]+z[55]);
assign {c[57],s[56]} = (x[56]+y[56]+z[56]);
assign {c[58],s[57]} = (x[57]+y[57]+z[57]);
assign {c[59],s[58]} = (x[58]+y[58]+z[58]);
assign {c[60],s[59]} = (x[59]+y[59]+z[59]);
assign {c[61],s[60]} = (x[60]+y[60]+z[60]);
assign {c[62],s[61]} = (x[61]+y[61]+z[61]);
assign {c[63],s[62]} = (x[62]+y[62]+z[62]);
assign {c[64],s[63]} = (x[63]+y[63]+z[63]);
assign {c[65],s[64]} = (x[64]+y[64]+z[64]);
assign {c[66],s[65]} = (x[65]+y[65]+z[65]);
assign {c[67],s[66]} = (x[66]+y[66]+z[66]);
assign {c[68],s[67]} = (x[67]+y[67]+z[67]);
assign {c[69],s[68]} = (x[68]+y[68]+z[68]);
assign {c[70],s[69]} = (x[69]+y[69]+z[69]);
assign {c[71],s[70]} = (x[70]+y[70]+z[70]);
assign {c[72],s[71]} = (x[71]+y[71]+z[71]);
assign {c[73],s[72]} = (x[72]+y[72]+z[72]);
assign {c[74],s[73]} = (x[73]+y[73]+z[73]);
assign {c[75],s[74]} = (x[74]+y[74]+z[74]);
assign {c[76],s[75]} = (x[75]+y[75]+z[75]);
assign {c[77],s[76]} = (x[76]+y[76]+z[76]);
assign {c[78],s[77]} = (x[77]+y[77]+z[77]);
assign {c[79],s[78]} = (x[78]+y[78]+z[78]);
assign {c[80],s[79]} = (x[79]+y[79]+z[79]);
assign {c[81],s[80]} = (x[80]+y[80]+z[80]);
assign {c[82],s[81]} = (x[81]+y[81]+z[81]);
assign {c[83],s[82]} = (x[82]+y[82]+z[82]);
assign {c[84],s[83]} = (x[83]+y[83]+z[83]);
assign {c[85],s[84]} = (x[84]+y[84]+z[84]);
assign {c[86],s[85]} = (x[85]+y[85]+z[85]);
assign {c[87],s[86]} = (x[86]+y[86]+z[86]);
assign {c[88],s[87]} = (x[87]+y[87]+z[87]);
assign {c[89],s[88]} = (x[88]+y[88]+z[88]);
assign {c[90],s[89]} = (x[89]+y[89]+z[89]);
assign {c[91],s[90]} = (x[90]+y[90]+z[90]);
assign {c[92],s[91]} = (x[91]+y[91]+z[91]);
assign {c[93],s[92]} = (x[92]+y[92]+z[92]);
assign {c[94],s[93]} = (x[93]+y[93]+z[93]);
assign {c[95],s[94]} = (x[94]+y[94]+z[94]);
assign {c[96],s[95]} = (x[95]+y[95]+z[95]);
assign {c[97],s[96]} = (x[96]+y[96]+z[96]);
assign {c[98],s[97]} = (x[97]+y[97]+z[97]);
assign {c[99],s[98]} = (x[98]+y[98]+z[98]);
assign {c[100],s[99]} = (x[99]+y[99]+z[99]);
assign {c[101],s[100]} = (x[100]+y[100]+z[100]);
assign {c[102],s[101]} = (x[101]+y[101]+z[101]);
assign {c[103],s[102]} = (x[102]+y[102]+z[102]);
assign {c[104],s[103]} = (x[103]+y[103]+z[103]);
assign {c[105],s[104]} = (x[104]+y[104]+z[104]);
assign {c[106],s[105]} = (x[105]+y[105]+z[105]);
assign {c[107],s[106]} = (x[106]+y[106]+z[106]);
assign {c[108],s[107]} = (x[107]+y[107]+z[107]);
assign {c[109],s[108]} = (x[108]+y[108]+z[108]);
assign {c[110],s[109]} = (x[109]+y[109]+z[109]);
assign {c[111],s[110]} = (x[110]+y[110]+z[110]);
assign {c[112],s[111]} = (x[111]+y[111]+z[111]);
assign {c[113],s[112]} = (x[112]+y[112]+z[112]);
assign {c[114],s[113]} = (x[113]+y[113]+z[113]);
assign {c[115],s[114]} = (x[114]+y[114]+z[114]);
assign {c[116],s[115]} = (x[115]+y[115]+z[115]);
assign {c[117],s[116]} = (x[116]+y[116]+z[116]);
assign {c[118],s[117]} = (x[117]+y[117]+z[117]);
assign {c[119],s[118]} = (x[118]+y[118]+z[118]);
assign {c[120],s[119]} = (x[119]+y[119]+z[119]);
assign {c[121],s[120]} = (x[120]+y[120]+z[120]);
assign {c[122],s[121]} = (x[121]+y[121]+z[121]);
assign {c[123],s[122]} = (x[122]+y[122]+z[122]);
assign {c[124],s[123]} = (x[123]+y[123]+z[123]);
assign {c[125],s[124]} = (x[124]+y[124]+z[124]);
assign {c[126],s[125]} = (x[125]+y[125]+z[125]);
assign {c[127],s[126]} = (x[126]+y[126]+z[126]);
assign {c[128],s[127]} = (x[127]+y[127]+z[127]);
assign {c[129],s[128]} = (x[128]+y[128]+z[128]);
assign {c[130],s[129]} = (x[129]+y[129]+z[129]);
assign {c[131],s[130]} = (x[130]+y[130]+z[130]);
assign {c[132],s[131]} = (x[131]+y[131]+z[131]);
assign {c[133],s[132]} = (x[132]+y[132]+z[132]);
assign {c[134],s[133]} = (x[133]+y[133]+z[133]);
assign {c[135],s[134]} = (x[134]+y[134]+z[134]);
assign {c[136],s[135]} = (x[135]+y[135]+z[135]);
assign {c[137],s[136]} = (x[136]+y[136]+z[136]);
assign {c[138],s[137]} = (x[137]+y[137]+z[137]);
assign {c[139],s[138]} = (x[138]+y[138]+z[138]);
assign {c[140],s[139]} = (x[139]+y[139]+z[139]);
assign {c[141],s[140]} = (x[140]+y[140]+z[140]);
assign {c[142],s[141]} = (x[141]+y[141]+z[141]);
assign {c[143],s[142]} = (x[142]+y[142]+z[142]);
assign {c[144],s[143]} = (x[143]+y[143]+z[143]);
assign {c[145],s[144]} = (x[144]+y[144]+z[144]);
assign {c[146],s[145]} = (x[145]+y[145]+z[145]);
assign {c[147],s[146]} = (x[146]+y[146]+z[146]);
assign {c[148],s[147]} = (x[147]+y[147]+z[147]);
assign {c[149],s[148]} = (x[148]+y[148]+z[148]);
assign {c[150],s[149]} = (x[149]+y[149]+z[149]);
assign {c[151],s[150]} = (x[150]+y[150]+z[150]);
assign {c[152],s[151]} = (x[151]+y[151]+z[151]);
assign {c[153],s[152]} = (x[152]+y[152]+z[152]);
assign {c[154],s[153]} = (x[153]+y[153]+z[153]);
assign {c[155],s[154]} = (x[154]+y[154]+z[154]);
assign {c[156],s[155]} = (x[155]+y[155]+z[155]);
assign {c[157],s[156]} = (x[156]+y[156]+z[156]);
assign {c[158],s[157]} = (x[157]+y[157]+z[157]);
assign {c[159],s[158]} = (x[158]+y[158]+z[158]);
assign {c[160],s[159]} = (x[159]+y[159]+z[159]);
assign {c[161],s[160]} = (x[160]+y[160]+z[160]);
assign {c[162],s[161]} = (x[161]+y[161]+z[161]);
assign {c[163],s[162]} = (x[162]+y[162]+z[162]);
assign {c[164],s[163]} = (x[163]+y[163]+z[163]);
assign {c[165],s[164]} = (x[164]+y[164]+z[164]);
assign {c[166],s[165]} = (x[165]+y[165]+z[165]);
assign {c[167],s[166]} = (x[166]+y[166]+z[166]);
assign {c[168],s[167]} = (x[167]+y[167]+z[167]);
assign {c[169],s[168]} = (x[168]+y[168]+z[168]);
assign {c[170],s[169]} = (x[169]+y[169]+z[169]);
assign {c[171],s[170]} = (x[170]+y[170]+z[170]);
assign {c[172],s[171]} = (x[171]+y[171]+z[171]);
assign {c[173],s[172]} = (x[172]+y[172]+z[172]);
assign {c[174],s[173]} = (x[173]+y[173]+z[173]);
assign {c[175],s[174]} = (x[174]+y[174]+z[174]);
assign {c[176],s[175]} = (x[175]+y[175]+z[175]);
assign {c[177],s[176]} = (x[176]+y[176]+z[176]);
assign {c[178],s[177]} = (x[177]+y[177]+z[177]);
assign {c[179],s[178]} = (x[178]+y[178]+z[178]);
assign {c[180],s[179]} = (x[179]+y[179]+z[179]);
assign {c[181],s[180]} = (x[180]+y[180]+z[180]);
assign {c[182],s[181]} = (x[181]+y[181]+z[181]);
assign {c[183],s[182]} = (x[182]+y[182]+z[182]);
assign {c[184],s[183]} = (x[183]+y[183]+z[183]);
assign {c[185],s[184]} = (x[184]+y[184]+z[184]);
assign {dummy,s[185]} = (x[185]+y[185]+z[185]);

endmodule
    