
module AND_matrix_1509x1509(
    input [1508:0] a,
    input [1508:0] b,
    output [4554161:0] c // lines are appended together
);
    
wire [1508:0] c_w_0;
wire [1508:0] c_w_1;
wire [1508:0] c_w_2;
wire [1508:0] c_w_3;
wire [1508:0] c_w_4;
wire [1508:0] c_w_5;
wire [1508:0] c_w_6;
wire [1508:0] c_w_7;
wire [1508:0] c_w_8;
wire [1508:0] c_w_9;
wire [1508:0] c_w_10;
wire [1508:0] c_w_11;
wire [1508:0] c_w_12;
wire [1508:0] c_w_13;
wire [1508:0] c_w_14;
wire [1508:0] c_w_15;
wire [1508:0] c_w_16;
wire [1508:0] c_w_17;
wire [1508:0] c_w_18;
wire [1508:0] c_w_19;
wire [1508:0] c_w_20;
wire [1508:0] c_w_21;
wire [1508:0] c_w_22;
wire [1508:0] c_w_23;
wire [1508:0] c_w_24;
wire [1508:0] c_w_25;
wire [1508:0] c_w_26;
wire [1508:0] c_w_27;
wire [1508:0] c_w_28;
wire [1508:0] c_w_29;
wire [1508:0] c_w_30;
wire [1508:0] c_w_31;
wire [1508:0] c_w_32;
wire [1508:0] c_w_33;
wire [1508:0] c_w_34;
wire [1508:0] c_w_35;
wire [1508:0] c_w_36;
wire [1508:0] c_w_37;
wire [1508:0] c_w_38;
wire [1508:0] c_w_39;
wire [1508:0] c_w_40;
wire [1508:0] c_w_41;
wire [1508:0] c_w_42;
wire [1508:0] c_w_43;
wire [1508:0] c_w_44;
wire [1508:0] c_w_45;
wire [1508:0] c_w_46;
wire [1508:0] c_w_47;
wire [1508:0] c_w_48;
wire [1508:0] c_w_49;
wire [1508:0] c_w_50;
wire [1508:0] c_w_51;
wire [1508:0] c_w_52;
wire [1508:0] c_w_53;
wire [1508:0] c_w_54;
wire [1508:0] c_w_55;
wire [1508:0] c_w_56;
wire [1508:0] c_w_57;
wire [1508:0] c_w_58;
wire [1508:0] c_w_59;
wire [1508:0] c_w_60;
wire [1508:0] c_w_61;
wire [1508:0] c_w_62;
wire [1508:0] c_w_63;
wire [1508:0] c_w_64;
wire [1508:0] c_w_65;
wire [1508:0] c_w_66;
wire [1508:0] c_w_67;
wire [1508:0] c_w_68;
wire [1508:0] c_w_69;
wire [1508:0] c_w_70;
wire [1508:0] c_w_71;
wire [1508:0] c_w_72;
wire [1508:0] c_w_73;
wire [1508:0] c_w_74;
wire [1508:0] c_w_75;
wire [1508:0] c_w_76;
wire [1508:0] c_w_77;
wire [1508:0] c_w_78;
wire [1508:0] c_w_79;
wire [1508:0] c_w_80;
wire [1508:0] c_w_81;
wire [1508:0] c_w_82;
wire [1508:0] c_w_83;
wire [1508:0] c_w_84;
wire [1508:0] c_w_85;
wire [1508:0] c_w_86;
wire [1508:0] c_w_87;
wire [1508:0] c_w_88;
wire [1508:0] c_w_89;
wire [1508:0] c_w_90;
wire [1508:0] c_w_91;
wire [1508:0] c_w_92;
wire [1508:0] c_w_93;
wire [1508:0] c_w_94;
wire [1508:0] c_w_95;
wire [1508:0] c_w_96;
wire [1508:0] c_w_97;
wire [1508:0] c_w_98;
wire [1508:0] c_w_99;
wire [1508:0] c_w_100;
wire [1508:0] c_w_101;
wire [1508:0] c_w_102;
wire [1508:0] c_w_103;
wire [1508:0] c_w_104;
wire [1508:0] c_w_105;
wire [1508:0] c_w_106;
wire [1508:0] c_w_107;
wire [1508:0] c_w_108;
wire [1508:0] c_w_109;
wire [1508:0] c_w_110;
wire [1508:0] c_w_111;
wire [1508:0] c_w_112;
wire [1508:0] c_w_113;
wire [1508:0] c_w_114;
wire [1508:0] c_w_115;
wire [1508:0] c_w_116;
wire [1508:0] c_w_117;
wire [1508:0] c_w_118;
wire [1508:0] c_w_119;
wire [1508:0] c_w_120;
wire [1508:0] c_w_121;
wire [1508:0] c_w_122;
wire [1508:0] c_w_123;
wire [1508:0] c_w_124;
wire [1508:0] c_w_125;
wire [1508:0] c_w_126;
wire [1508:0] c_w_127;
wire [1508:0] c_w_128;
wire [1508:0] c_w_129;
wire [1508:0] c_w_130;
wire [1508:0] c_w_131;
wire [1508:0] c_w_132;
wire [1508:0] c_w_133;
wire [1508:0] c_w_134;
wire [1508:0] c_w_135;
wire [1508:0] c_w_136;
wire [1508:0] c_w_137;
wire [1508:0] c_w_138;
wire [1508:0] c_w_139;
wire [1508:0] c_w_140;
wire [1508:0] c_w_141;
wire [1508:0] c_w_142;
wire [1508:0] c_w_143;
wire [1508:0] c_w_144;
wire [1508:0] c_w_145;
wire [1508:0] c_w_146;
wire [1508:0] c_w_147;
wire [1508:0] c_w_148;
wire [1508:0] c_w_149;
wire [1508:0] c_w_150;
wire [1508:0] c_w_151;
wire [1508:0] c_w_152;
wire [1508:0] c_w_153;
wire [1508:0] c_w_154;
wire [1508:0] c_w_155;
wire [1508:0] c_w_156;
wire [1508:0] c_w_157;
wire [1508:0] c_w_158;
wire [1508:0] c_w_159;
wire [1508:0] c_w_160;
wire [1508:0] c_w_161;
wire [1508:0] c_w_162;
wire [1508:0] c_w_163;
wire [1508:0] c_w_164;
wire [1508:0] c_w_165;
wire [1508:0] c_w_166;
wire [1508:0] c_w_167;
wire [1508:0] c_w_168;
wire [1508:0] c_w_169;
wire [1508:0] c_w_170;
wire [1508:0] c_w_171;
wire [1508:0] c_w_172;
wire [1508:0] c_w_173;
wire [1508:0] c_w_174;
wire [1508:0] c_w_175;
wire [1508:0] c_w_176;
wire [1508:0] c_w_177;
wire [1508:0] c_w_178;
wire [1508:0] c_w_179;
wire [1508:0] c_w_180;
wire [1508:0] c_w_181;
wire [1508:0] c_w_182;
wire [1508:0] c_w_183;
wire [1508:0] c_w_184;
wire [1508:0] c_w_185;
wire [1508:0] c_w_186;
wire [1508:0] c_w_187;
wire [1508:0] c_w_188;
wire [1508:0] c_w_189;
wire [1508:0] c_w_190;
wire [1508:0] c_w_191;
wire [1508:0] c_w_192;
wire [1508:0] c_w_193;
wire [1508:0] c_w_194;
wire [1508:0] c_w_195;
wire [1508:0] c_w_196;
wire [1508:0] c_w_197;
wire [1508:0] c_w_198;
wire [1508:0] c_w_199;
wire [1508:0] c_w_200;
wire [1508:0] c_w_201;
wire [1508:0] c_w_202;
wire [1508:0] c_w_203;
wire [1508:0] c_w_204;
wire [1508:0] c_w_205;
wire [1508:0] c_w_206;
wire [1508:0] c_w_207;
wire [1508:0] c_w_208;
wire [1508:0] c_w_209;
wire [1508:0] c_w_210;
wire [1508:0] c_w_211;
wire [1508:0] c_w_212;
wire [1508:0] c_w_213;
wire [1508:0] c_w_214;
wire [1508:0] c_w_215;
wire [1508:0] c_w_216;
wire [1508:0] c_w_217;
wire [1508:0] c_w_218;
wire [1508:0] c_w_219;
wire [1508:0] c_w_220;
wire [1508:0] c_w_221;
wire [1508:0] c_w_222;
wire [1508:0] c_w_223;
wire [1508:0] c_w_224;
wire [1508:0] c_w_225;
wire [1508:0] c_w_226;
wire [1508:0] c_w_227;
wire [1508:0] c_w_228;
wire [1508:0] c_w_229;
wire [1508:0] c_w_230;
wire [1508:0] c_w_231;
wire [1508:0] c_w_232;
wire [1508:0] c_w_233;
wire [1508:0] c_w_234;
wire [1508:0] c_w_235;
wire [1508:0] c_w_236;
wire [1508:0] c_w_237;
wire [1508:0] c_w_238;
wire [1508:0] c_w_239;
wire [1508:0] c_w_240;
wire [1508:0] c_w_241;
wire [1508:0] c_w_242;
wire [1508:0] c_w_243;
wire [1508:0] c_w_244;
wire [1508:0] c_w_245;
wire [1508:0] c_w_246;
wire [1508:0] c_w_247;
wire [1508:0] c_w_248;
wire [1508:0] c_w_249;
wire [1508:0] c_w_250;
wire [1508:0] c_w_251;
wire [1508:0] c_w_252;
wire [1508:0] c_w_253;
wire [1508:0] c_w_254;
wire [1508:0] c_w_255;
wire [1508:0] c_w_256;
wire [1508:0] c_w_257;
wire [1508:0] c_w_258;
wire [1508:0] c_w_259;
wire [1508:0] c_w_260;
wire [1508:0] c_w_261;
wire [1508:0] c_w_262;
wire [1508:0] c_w_263;
wire [1508:0] c_w_264;
wire [1508:0] c_w_265;
wire [1508:0] c_w_266;
wire [1508:0] c_w_267;
wire [1508:0] c_w_268;
wire [1508:0] c_w_269;
wire [1508:0] c_w_270;
wire [1508:0] c_w_271;
wire [1508:0] c_w_272;
wire [1508:0] c_w_273;
wire [1508:0] c_w_274;
wire [1508:0] c_w_275;
wire [1508:0] c_w_276;
wire [1508:0] c_w_277;
wire [1508:0] c_w_278;
wire [1508:0] c_w_279;
wire [1508:0] c_w_280;
wire [1508:0] c_w_281;
wire [1508:0] c_w_282;
wire [1508:0] c_w_283;
wire [1508:0] c_w_284;
wire [1508:0] c_w_285;
wire [1508:0] c_w_286;
wire [1508:0] c_w_287;
wire [1508:0] c_w_288;
wire [1508:0] c_w_289;
wire [1508:0] c_w_290;
wire [1508:0] c_w_291;
wire [1508:0] c_w_292;
wire [1508:0] c_w_293;
wire [1508:0] c_w_294;
wire [1508:0] c_w_295;
wire [1508:0] c_w_296;
wire [1508:0] c_w_297;
wire [1508:0] c_w_298;
wire [1508:0] c_w_299;
wire [1508:0] c_w_300;
wire [1508:0] c_w_301;
wire [1508:0] c_w_302;
wire [1508:0] c_w_303;
wire [1508:0] c_w_304;
wire [1508:0] c_w_305;
wire [1508:0] c_w_306;
wire [1508:0] c_w_307;
wire [1508:0] c_w_308;
wire [1508:0] c_w_309;
wire [1508:0] c_w_310;
wire [1508:0] c_w_311;
wire [1508:0] c_w_312;
wire [1508:0] c_w_313;
wire [1508:0] c_w_314;
wire [1508:0] c_w_315;
wire [1508:0] c_w_316;
wire [1508:0] c_w_317;
wire [1508:0] c_w_318;
wire [1508:0] c_w_319;
wire [1508:0] c_w_320;
wire [1508:0] c_w_321;
wire [1508:0] c_w_322;
wire [1508:0] c_w_323;
wire [1508:0] c_w_324;
wire [1508:0] c_w_325;
wire [1508:0] c_w_326;
wire [1508:0] c_w_327;
wire [1508:0] c_w_328;
wire [1508:0] c_w_329;
wire [1508:0] c_w_330;
wire [1508:0] c_w_331;
wire [1508:0] c_w_332;
wire [1508:0] c_w_333;
wire [1508:0] c_w_334;
wire [1508:0] c_w_335;
wire [1508:0] c_w_336;
wire [1508:0] c_w_337;
wire [1508:0] c_w_338;
wire [1508:0] c_w_339;
wire [1508:0] c_w_340;
wire [1508:0] c_w_341;
wire [1508:0] c_w_342;
wire [1508:0] c_w_343;
wire [1508:0] c_w_344;
wire [1508:0] c_w_345;
wire [1508:0] c_w_346;
wire [1508:0] c_w_347;
wire [1508:0] c_w_348;
wire [1508:0] c_w_349;
wire [1508:0] c_w_350;
wire [1508:0] c_w_351;
wire [1508:0] c_w_352;
wire [1508:0] c_w_353;
wire [1508:0] c_w_354;
wire [1508:0] c_w_355;
wire [1508:0] c_w_356;
wire [1508:0] c_w_357;
wire [1508:0] c_w_358;
wire [1508:0] c_w_359;
wire [1508:0] c_w_360;
wire [1508:0] c_w_361;
wire [1508:0] c_w_362;
wire [1508:0] c_w_363;
wire [1508:0] c_w_364;
wire [1508:0] c_w_365;
wire [1508:0] c_w_366;
wire [1508:0] c_w_367;
wire [1508:0] c_w_368;
wire [1508:0] c_w_369;
wire [1508:0] c_w_370;
wire [1508:0] c_w_371;
wire [1508:0] c_w_372;
wire [1508:0] c_w_373;
wire [1508:0] c_w_374;
wire [1508:0] c_w_375;
wire [1508:0] c_w_376;
wire [1508:0] c_w_377;
wire [1508:0] c_w_378;
wire [1508:0] c_w_379;
wire [1508:0] c_w_380;
wire [1508:0] c_w_381;
wire [1508:0] c_w_382;
wire [1508:0] c_w_383;
wire [1508:0] c_w_384;
wire [1508:0] c_w_385;
wire [1508:0] c_w_386;
wire [1508:0] c_w_387;
wire [1508:0] c_w_388;
wire [1508:0] c_w_389;
wire [1508:0] c_w_390;
wire [1508:0] c_w_391;
wire [1508:0] c_w_392;
wire [1508:0] c_w_393;
wire [1508:0] c_w_394;
wire [1508:0] c_w_395;
wire [1508:0] c_w_396;
wire [1508:0] c_w_397;
wire [1508:0] c_w_398;
wire [1508:0] c_w_399;
wire [1508:0] c_w_400;
wire [1508:0] c_w_401;
wire [1508:0] c_w_402;
wire [1508:0] c_w_403;
wire [1508:0] c_w_404;
wire [1508:0] c_w_405;
wire [1508:0] c_w_406;
wire [1508:0] c_w_407;
wire [1508:0] c_w_408;
wire [1508:0] c_w_409;
wire [1508:0] c_w_410;
wire [1508:0] c_w_411;
wire [1508:0] c_w_412;
wire [1508:0] c_w_413;
wire [1508:0] c_w_414;
wire [1508:0] c_w_415;
wire [1508:0] c_w_416;
wire [1508:0] c_w_417;
wire [1508:0] c_w_418;
wire [1508:0] c_w_419;
wire [1508:0] c_w_420;
wire [1508:0] c_w_421;
wire [1508:0] c_w_422;
wire [1508:0] c_w_423;
wire [1508:0] c_w_424;
wire [1508:0] c_w_425;
wire [1508:0] c_w_426;
wire [1508:0] c_w_427;
wire [1508:0] c_w_428;
wire [1508:0] c_w_429;
wire [1508:0] c_w_430;
wire [1508:0] c_w_431;
wire [1508:0] c_w_432;
wire [1508:0] c_w_433;
wire [1508:0] c_w_434;
wire [1508:0] c_w_435;
wire [1508:0] c_w_436;
wire [1508:0] c_w_437;
wire [1508:0] c_w_438;
wire [1508:0] c_w_439;
wire [1508:0] c_w_440;
wire [1508:0] c_w_441;
wire [1508:0] c_w_442;
wire [1508:0] c_w_443;
wire [1508:0] c_w_444;
wire [1508:0] c_w_445;
wire [1508:0] c_w_446;
wire [1508:0] c_w_447;
wire [1508:0] c_w_448;
wire [1508:0] c_w_449;
wire [1508:0] c_w_450;
wire [1508:0] c_w_451;
wire [1508:0] c_w_452;
wire [1508:0] c_w_453;
wire [1508:0] c_w_454;
wire [1508:0] c_w_455;
wire [1508:0] c_w_456;
wire [1508:0] c_w_457;
wire [1508:0] c_w_458;
wire [1508:0] c_w_459;
wire [1508:0] c_w_460;
wire [1508:0] c_w_461;
wire [1508:0] c_w_462;
wire [1508:0] c_w_463;
wire [1508:0] c_w_464;
wire [1508:0] c_w_465;
wire [1508:0] c_w_466;
wire [1508:0] c_w_467;
wire [1508:0] c_w_468;
wire [1508:0] c_w_469;
wire [1508:0] c_w_470;
wire [1508:0] c_w_471;
wire [1508:0] c_w_472;
wire [1508:0] c_w_473;
wire [1508:0] c_w_474;
wire [1508:0] c_w_475;
wire [1508:0] c_w_476;
wire [1508:0] c_w_477;
wire [1508:0] c_w_478;
wire [1508:0] c_w_479;
wire [1508:0] c_w_480;
wire [1508:0] c_w_481;
wire [1508:0] c_w_482;
wire [1508:0] c_w_483;
wire [1508:0] c_w_484;
wire [1508:0] c_w_485;
wire [1508:0] c_w_486;
wire [1508:0] c_w_487;
wire [1508:0] c_w_488;
wire [1508:0] c_w_489;
wire [1508:0] c_w_490;
wire [1508:0] c_w_491;
wire [1508:0] c_w_492;
wire [1508:0] c_w_493;
wire [1508:0] c_w_494;
wire [1508:0] c_w_495;
wire [1508:0] c_w_496;
wire [1508:0] c_w_497;
wire [1508:0] c_w_498;
wire [1508:0] c_w_499;
wire [1508:0] c_w_500;
wire [1508:0] c_w_501;
wire [1508:0] c_w_502;
wire [1508:0] c_w_503;
wire [1508:0] c_w_504;
wire [1508:0] c_w_505;
wire [1508:0] c_w_506;
wire [1508:0] c_w_507;
wire [1508:0] c_w_508;
wire [1508:0] c_w_509;
wire [1508:0] c_w_510;
wire [1508:0] c_w_511;
wire [1508:0] c_w_512;
wire [1508:0] c_w_513;
wire [1508:0] c_w_514;
wire [1508:0] c_w_515;
wire [1508:0] c_w_516;
wire [1508:0] c_w_517;
wire [1508:0] c_w_518;
wire [1508:0] c_w_519;
wire [1508:0] c_w_520;
wire [1508:0] c_w_521;
wire [1508:0] c_w_522;
wire [1508:0] c_w_523;
wire [1508:0] c_w_524;
wire [1508:0] c_w_525;
wire [1508:0] c_w_526;
wire [1508:0] c_w_527;
wire [1508:0] c_w_528;
wire [1508:0] c_w_529;
wire [1508:0] c_w_530;
wire [1508:0] c_w_531;
wire [1508:0] c_w_532;
wire [1508:0] c_w_533;
wire [1508:0] c_w_534;
wire [1508:0] c_w_535;
wire [1508:0] c_w_536;
wire [1508:0] c_w_537;
wire [1508:0] c_w_538;
wire [1508:0] c_w_539;
wire [1508:0] c_w_540;
wire [1508:0] c_w_541;
wire [1508:0] c_w_542;
wire [1508:0] c_w_543;
wire [1508:0] c_w_544;
wire [1508:0] c_w_545;
wire [1508:0] c_w_546;
wire [1508:0] c_w_547;
wire [1508:0] c_w_548;
wire [1508:0] c_w_549;
wire [1508:0] c_w_550;
wire [1508:0] c_w_551;
wire [1508:0] c_w_552;
wire [1508:0] c_w_553;
wire [1508:0] c_w_554;
wire [1508:0] c_w_555;
wire [1508:0] c_w_556;
wire [1508:0] c_w_557;
wire [1508:0] c_w_558;
wire [1508:0] c_w_559;
wire [1508:0] c_w_560;
wire [1508:0] c_w_561;
wire [1508:0] c_w_562;
wire [1508:0] c_w_563;
wire [1508:0] c_w_564;
wire [1508:0] c_w_565;
wire [1508:0] c_w_566;
wire [1508:0] c_w_567;
wire [1508:0] c_w_568;
wire [1508:0] c_w_569;
wire [1508:0] c_w_570;
wire [1508:0] c_w_571;
wire [1508:0] c_w_572;
wire [1508:0] c_w_573;
wire [1508:0] c_w_574;
wire [1508:0] c_w_575;
wire [1508:0] c_w_576;
wire [1508:0] c_w_577;
wire [1508:0] c_w_578;
wire [1508:0] c_w_579;
wire [1508:0] c_w_580;
wire [1508:0] c_w_581;
wire [1508:0] c_w_582;
wire [1508:0] c_w_583;
wire [1508:0] c_w_584;
wire [1508:0] c_w_585;
wire [1508:0] c_w_586;
wire [1508:0] c_w_587;
wire [1508:0] c_w_588;
wire [1508:0] c_w_589;
wire [1508:0] c_w_590;
wire [1508:0] c_w_591;
wire [1508:0] c_w_592;
wire [1508:0] c_w_593;
wire [1508:0] c_w_594;
wire [1508:0] c_w_595;
wire [1508:0] c_w_596;
wire [1508:0] c_w_597;
wire [1508:0] c_w_598;
wire [1508:0] c_w_599;
wire [1508:0] c_w_600;
wire [1508:0] c_w_601;
wire [1508:0] c_w_602;
wire [1508:0] c_w_603;
wire [1508:0] c_w_604;
wire [1508:0] c_w_605;
wire [1508:0] c_w_606;
wire [1508:0] c_w_607;
wire [1508:0] c_w_608;
wire [1508:0] c_w_609;
wire [1508:0] c_w_610;
wire [1508:0] c_w_611;
wire [1508:0] c_w_612;
wire [1508:0] c_w_613;
wire [1508:0] c_w_614;
wire [1508:0] c_w_615;
wire [1508:0] c_w_616;
wire [1508:0] c_w_617;
wire [1508:0] c_w_618;
wire [1508:0] c_w_619;
wire [1508:0] c_w_620;
wire [1508:0] c_w_621;
wire [1508:0] c_w_622;
wire [1508:0] c_w_623;
wire [1508:0] c_w_624;
wire [1508:0] c_w_625;
wire [1508:0] c_w_626;
wire [1508:0] c_w_627;
wire [1508:0] c_w_628;
wire [1508:0] c_w_629;
wire [1508:0] c_w_630;
wire [1508:0] c_w_631;
wire [1508:0] c_w_632;
wire [1508:0] c_w_633;
wire [1508:0] c_w_634;
wire [1508:0] c_w_635;
wire [1508:0] c_w_636;
wire [1508:0] c_w_637;
wire [1508:0] c_w_638;
wire [1508:0] c_w_639;
wire [1508:0] c_w_640;
wire [1508:0] c_w_641;
wire [1508:0] c_w_642;
wire [1508:0] c_w_643;
wire [1508:0] c_w_644;
wire [1508:0] c_w_645;
wire [1508:0] c_w_646;
wire [1508:0] c_w_647;
wire [1508:0] c_w_648;
wire [1508:0] c_w_649;
wire [1508:0] c_w_650;
wire [1508:0] c_w_651;
wire [1508:0] c_w_652;
wire [1508:0] c_w_653;
wire [1508:0] c_w_654;
wire [1508:0] c_w_655;
wire [1508:0] c_w_656;
wire [1508:0] c_w_657;
wire [1508:0] c_w_658;
wire [1508:0] c_w_659;
wire [1508:0] c_w_660;
wire [1508:0] c_w_661;
wire [1508:0] c_w_662;
wire [1508:0] c_w_663;
wire [1508:0] c_w_664;
wire [1508:0] c_w_665;
wire [1508:0] c_w_666;
wire [1508:0] c_w_667;
wire [1508:0] c_w_668;
wire [1508:0] c_w_669;
wire [1508:0] c_w_670;
wire [1508:0] c_w_671;
wire [1508:0] c_w_672;
wire [1508:0] c_w_673;
wire [1508:0] c_w_674;
wire [1508:0] c_w_675;
wire [1508:0] c_w_676;
wire [1508:0] c_w_677;
wire [1508:0] c_w_678;
wire [1508:0] c_w_679;
wire [1508:0] c_w_680;
wire [1508:0] c_w_681;
wire [1508:0] c_w_682;
wire [1508:0] c_w_683;
wire [1508:0] c_w_684;
wire [1508:0] c_w_685;
wire [1508:0] c_w_686;
wire [1508:0] c_w_687;
wire [1508:0] c_w_688;
wire [1508:0] c_w_689;
wire [1508:0] c_w_690;
wire [1508:0] c_w_691;
wire [1508:0] c_w_692;
wire [1508:0] c_w_693;
wire [1508:0] c_w_694;
wire [1508:0] c_w_695;
wire [1508:0] c_w_696;
wire [1508:0] c_w_697;
wire [1508:0] c_w_698;
wire [1508:0] c_w_699;
wire [1508:0] c_w_700;
wire [1508:0] c_w_701;
wire [1508:0] c_w_702;
wire [1508:0] c_w_703;
wire [1508:0] c_w_704;
wire [1508:0] c_w_705;
wire [1508:0] c_w_706;
wire [1508:0] c_w_707;
wire [1508:0] c_w_708;
wire [1508:0] c_w_709;
wire [1508:0] c_w_710;
wire [1508:0] c_w_711;
wire [1508:0] c_w_712;
wire [1508:0] c_w_713;
wire [1508:0] c_w_714;
wire [1508:0] c_w_715;
wire [1508:0] c_w_716;
wire [1508:0] c_w_717;
wire [1508:0] c_w_718;
wire [1508:0] c_w_719;
wire [1508:0] c_w_720;
wire [1508:0] c_w_721;
wire [1508:0] c_w_722;
wire [1508:0] c_w_723;
wire [1508:0] c_w_724;
wire [1508:0] c_w_725;
wire [1508:0] c_w_726;
wire [1508:0] c_w_727;
wire [1508:0] c_w_728;
wire [1508:0] c_w_729;
wire [1508:0] c_w_730;
wire [1508:0] c_w_731;
wire [1508:0] c_w_732;
wire [1508:0] c_w_733;
wire [1508:0] c_w_734;
wire [1508:0] c_w_735;
wire [1508:0] c_w_736;
wire [1508:0] c_w_737;
wire [1508:0] c_w_738;
wire [1508:0] c_w_739;
wire [1508:0] c_w_740;
wire [1508:0] c_w_741;
wire [1508:0] c_w_742;
wire [1508:0] c_w_743;
wire [1508:0] c_w_744;
wire [1508:0] c_w_745;
wire [1508:0] c_w_746;
wire [1508:0] c_w_747;
wire [1508:0] c_w_748;
wire [1508:0] c_w_749;
wire [1508:0] c_w_750;
wire [1508:0] c_w_751;
wire [1508:0] c_w_752;
wire [1508:0] c_w_753;
wire [1508:0] c_w_754;
wire [1508:0] c_w_755;
wire [1508:0] c_w_756;
wire [1508:0] c_w_757;
wire [1508:0] c_w_758;
wire [1508:0] c_w_759;
wire [1508:0] c_w_760;
wire [1508:0] c_w_761;
wire [1508:0] c_w_762;
wire [1508:0] c_w_763;
wire [1508:0] c_w_764;
wire [1508:0] c_w_765;
wire [1508:0] c_w_766;
wire [1508:0] c_w_767;
wire [1508:0] c_w_768;
wire [1508:0] c_w_769;
wire [1508:0] c_w_770;
wire [1508:0] c_w_771;
wire [1508:0] c_w_772;
wire [1508:0] c_w_773;
wire [1508:0] c_w_774;
wire [1508:0] c_w_775;
wire [1508:0] c_w_776;
wire [1508:0] c_w_777;
wire [1508:0] c_w_778;
wire [1508:0] c_w_779;
wire [1508:0] c_w_780;
wire [1508:0] c_w_781;
wire [1508:0] c_w_782;
wire [1508:0] c_w_783;
wire [1508:0] c_w_784;
wire [1508:0] c_w_785;
wire [1508:0] c_w_786;
wire [1508:0] c_w_787;
wire [1508:0] c_w_788;
wire [1508:0] c_w_789;
wire [1508:0] c_w_790;
wire [1508:0] c_w_791;
wire [1508:0] c_w_792;
wire [1508:0] c_w_793;
wire [1508:0] c_w_794;
wire [1508:0] c_w_795;
wire [1508:0] c_w_796;
wire [1508:0] c_w_797;
wire [1508:0] c_w_798;
wire [1508:0] c_w_799;
wire [1508:0] c_w_800;
wire [1508:0] c_w_801;
wire [1508:0] c_w_802;
wire [1508:0] c_w_803;
wire [1508:0] c_w_804;
wire [1508:0] c_w_805;
wire [1508:0] c_w_806;
wire [1508:0] c_w_807;
wire [1508:0] c_w_808;
wire [1508:0] c_w_809;
wire [1508:0] c_w_810;
wire [1508:0] c_w_811;
wire [1508:0] c_w_812;
wire [1508:0] c_w_813;
wire [1508:0] c_w_814;
wire [1508:0] c_w_815;
wire [1508:0] c_w_816;
wire [1508:0] c_w_817;
wire [1508:0] c_w_818;
wire [1508:0] c_w_819;
wire [1508:0] c_w_820;
wire [1508:0] c_w_821;
wire [1508:0] c_w_822;
wire [1508:0] c_w_823;
wire [1508:0] c_w_824;
wire [1508:0] c_w_825;
wire [1508:0] c_w_826;
wire [1508:0] c_w_827;
wire [1508:0] c_w_828;
wire [1508:0] c_w_829;
wire [1508:0] c_w_830;
wire [1508:0] c_w_831;
wire [1508:0] c_w_832;
wire [1508:0] c_w_833;
wire [1508:0] c_w_834;
wire [1508:0] c_w_835;
wire [1508:0] c_w_836;
wire [1508:0] c_w_837;
wire [1508:0] c_w_838;
wire [1508:0] c_w_839;
wire [1508:0] c_w_840;
wire [1508:0] c_w_841;
wire [1508:0] c_w_842;
wire [1508:0] c_w_843;
wire [1508:0] c_w_844;
wire [1508:0] c_w_845;
wire [1508:0] c_w_846;
wire [1508:0] c_w_847;
wire [1508:0] c_w_848;
wire [1508:0] c_w_849;
wire [1508:0] c_w_850;
wire [1508:0] c_w_851;
wire [1508:0] c_w_852;
wire [1508:0] c_w_853;
wire [1508:0] c_w_854;
wire [1508:0] c_w_855;
wire [1508:0] c_w_856;
wire [1508:0] c_w_857;
wire [1508:0] c_w_858;
wire [1508:0] c_w_859;
wire [1508:0] c_w_860;
wire [1508:0] c_w_861;
wire [1508:0] c_w_862;
wire [1508:0] c_w_863;
wire [1508:0] c_w_864;
wire [1508:0] c_w_865;
wire [1508:0] c_w_866;
wire [1508:0] c_w_867;
wire [1508:0] c_w_868;
wire [1508:0] c_w_869;
wire [1508:0] c_w_870;
wire [1508:0] c_w_871;
wire [1508:0] c_w_872;
wire [1508:0] c_w_873;
wire [1508:0] c_w_874;
wire [1508:0] c_w_875;
wire [1508:0] c_w_876;
wire [1508:0] c_w_877;
wire [1508:0] c_w_878;
wire [1508:0] c_w_879;
wire [1508:0] c_w_880;
wire [1508:0] c_w_881;
wire [1508:0] c_w_882;
wire [1508:0] c_w_883;
wire [1508:0] c_w_884;
wire [1508:0] c_w_885;
wire [1508:0] c_w_886;
wire [1508:0] c_w_887;
wire [1508:0] c_w_888;
wire [1508:0] c_w_889;
wire [1508:0] c_w_890;
wire [1508:0] c_w_891;
wire [1508:0] c_w_892;
wire [1508:0] c_w_893;
wire [1508:0] c_w_894;
wire [1508:0] c_w_895;
wire [1508:0] c_w_896;
wire [1508:0] c_w_897;
wire [1508:0] c_w_898;
wire [1508:0] c_w_899;
wire [1508:0] c_w_900;
wire [1508:0] c_w_901;
wire [1508:0] c_w_902;
wire [1508:0] c_w_903;
wire [1508:0] c_w_904;
wire [1508:0] c_w_905;
wire [1508:0] c_w_906;
wire [1508:0] c_w_907;
wire [1508:0] c_w_908;
wire [1508:0] c_w_909;
wire [1508:0] c_w_910;
wire [1508:0] c_w_911;
wire [1508:0] c_w_912;
wire [1508:0] c_w_913;
wire [1508:0] c_w_914;
wire [1508:0] c_w_915;
wire [1508:0] c_w_916;
wire [1508:0] c_w_917;
wire [1508:0] c_w_918;
wire [1508:0] c_w_919;
wire [1508:0] c_w_920;
wire [1508:0] c_w_921;
wire [1508:0] c_w_922;
wire [1508:0] c_w_923;
wire [1508:0] c_w_924;
wire [1508:0] c_w_925;
wire [1508:0] c_w_926;
wire [1508:0] c_w_927;
wire [1508:0] c_w_928;
wire [1508:0] c_w_929;
wire [1508:0] c_w_930;
wire [1508:0] c_w_931;
wire [1508:0] c_w_932;
wire [1508:0] c_w_933;
wire [1508:0] c_w_934;
wire [1508:0] c_w_935;
wire [1508:0] c_w_936;
wire [1508:0] c_w_937;
wire [1508:0] c_w_938;
wire [1508:0] c_w_939;
wire [1508:0] c_w_940;
wire [1508:0] c_w_941;
wire [1508:0] c_w_942;
wire [1508:0] c_w_943;
wire [1508:0] c_w_944;
wire [1508:0] c_w_945;
wire [1508:0] c_w_946;
wire [1508:0] c_w_947;
wire [1508:0] c_w_948;
wire [1508:0] c_w_949;
wire [1508:0] c_w_950;
wire [1508:0] c_w_951;
wire [1508:0] c_w_952;
wire [1508:0] c_w_953;
wire [1508:0] c_w_954;
wire [1508:0] c_w_955;
wire [1508:0] c_w_956;
wire [1508:0] c_w_957;
wire [1508:0] c_w_958;
wire [1508:0] c_w_959;
wire [1508:0] c_w_960;
wire [1508:0] c_w_961;
wire [1508:0] c_w_962;
wire [1508:0] c_w_963;
wire [1508:0] c_w_964;
wire [1508:0] c_w_965;
wire [1508:0] c_w_966;
wire [1508:0] c_w_967;
wire [1508:0] c_w_968;
wire [1508:0] c_w_969;
wire [1508:0] c_w_970;
wire [1508:0] c_w_971;
wire [1508:0] c_w_972;
wire [1508:0] c_w_973;
wire [1508:0] c_w_974;
wire [1508:0] c_w_975;
wire [1508:0] c_w_976;
wire [1508:0] c_w_977;
wire [1508:0] c_w_978;
wire [1508:0] c_w_979;
wire [1508:0] c_w_980;
wire [1508:0] c_w_981;
wire [1508:0] c_w_982;
wire [1508:0] c_w_983;
wire [1508:0] c_w_984;
wire [1508:0] c_w_985;
wire [1508:0] c_w_986;
wire [1508:0] c_w_987;
wire [1508:0] c_w_988;
wire [1508:0] c_w_989;
wire [1508:0] c_w_990;
wire [1508:0] c_w_991;
wire [1508:0] c_w_992;
wire [1508:0] c_w_993;
wire [1508:0] c_w_994;
wire [1508:0] c_w_995;
wire [1508:0] c_w_996;
wire [1508:0] c_w_997;
wire [1508:0] c_w_998;
wire [1508:0] c_w_999;
wire [1508:0] c_w_1000;
wire [1508:0] c_w_1001;
wire [1508:0] c_w_1002;
wire [1508:0] c_w_1003;
wire [1508:0] c_w_1004;
wire [1508:0] c_w_1005;
wire [1508:0] c_w_1006;
wire [1508:0] c_w_1007;
wire [1508:0] c_w_1008;
wire [1508:0] c_w_1009;
wire [1508:0] c_w_1010;
wire [1508:0] c_w_1011;
wire [1508:0] c_w_1012;
wire [1508:0] c_w_1013;
wire [1508:0] c_w_1014;
wire [1508:0] c_w_1015;
wire [1508:0] c_w_1016;
wire [1508:0] c_w_1017;
wire [1508:0] c_w_1018;
wire [1508:0] c_w_1019;
wire [1508:0] c_w_1020;
wire [1508:0] c_w_1021;
wire [1508:0] c_w_1022;
wire [1508:0] c_w_1023;
wire [1508:0] c_w_1024;
wire [1508:0] c_w_1025;
wire [1508:0] c_w_1026;
wire [1508:0] c_w_1027;
wire [1508:0] c_w_1028;
wire [1508:0] c_w_1029;
wire [1508:0] c_w_1030;
wire [1508:0] c_w_1031;
wire [1508:0] c_w_1032;
wire [1508:0] c_w_1033;
wire [1508:0] c_w_1034;
wire [1508:0] c_w_1035;
wire [1508:0] c_w_1036;
wire [1508:0] c_w_1037;
wire [1508:0] c_w_1038;
wire [1508:0] c_w_1039;
wire [1508:0] c_w_1040;
wire [1508:0] c_w_1041;
wire [1508:0] c_w_1042;
wire [1508:0] c_w_1043;
wire [1508:0] c_w_1044;
wire [1508:0] c_w_1045;
wire [1508:0] c_w_1046;
wire [1508:0] c_w_1047;
wire [1508:0] c_w_1048;
wire [1508:0] c_w_1049;
wire [1508:0] c_w_1050;
wire [1508:0] c_w_1051;
wire [1508:0] c_w_1052;
wire [1508:0] c_w_1053;
wire [1508:0] c_w_1054;
wire [1508:0] c_w_1055;
wire [1508:0] c_w_1056;
wire [1508:0] c_w_1057;
wire [1508:0] c_w_1058;
wire [1508:0] c_w_1059;
wire [1508:0] c_w_1060;
wire [1508:0] c_w_1061;
wire [1508:0] c_w_1062;
wire [1508:0] c_w_1063;
wire [1508:0] c_w_1064;
wire [1508:0] c_w_1065;
wire [1508:0] c_w_1066;
wire [1508:0] c_w_1067;
wire [1508:0] c_w_1068;
wire [1508:0] c_w_1069;
wire [1508:0] c_w_1070;
wire [1508:0] c_w_1071;
wire [1508:0] c_w_1072;
wire [1508:0] c_w_1073;
wire [1508:0] c_w_1074;
wire [1508:0] c_w_1075;
wire [1508:0] c_w_1076;
wire [1508:0] c_w_1077;
wire [1508:0] c_w_1078;
wire [1508:0] c_w_1079;
wire [1508:0] c_w_1080;
wire [1508:0] c_w_1081;
wire [1508:0] c_w_1082;
wire [1508:0] c_w_1083;
wire [1508:0] c_w_1084;
wire [1508:0] c_w_1085;
wire [1508:0] c_w_1086;
wire [1508:0] c_w_1087;
wire [1508:0] c_w_1088;
wire [1508:0] c_w_1089;
wire [1508:0] c_w_1090;
wire [1508:0] c_w_1091;
wire [1508:0] c_w_1092;
wire [1508:0] c_w_1093;
wire [1508:0] c_w_1094;
wire [1508:0] c_w_1095;
wire [1508:0] c_w_1096;
wire [1508:0] c_w_1097;
wire [1508:0] c_w_1098;
wire [1508:0] c_w_1099;
wire [1508:0] c_w_1100;
wire [1508:0] c_w_1101;
wire [1508:0] c_w_1102;
wire [1508:0] c_w_1103;
wire [1508:0] c_w_1104;
wire [1508:0] c_w_1105;
wire [1508:0] c_w_1106;
wire [1508:0] c_w_1107;
wire [1508:0] c_w_1108;
wire [1508:0] c_w_1109;
wire [1508:0] c_w_1110;
wire [1508:0] c_w_1111;
wire [1508:0] c_w_1112;
wire [1508:0] c_w_1113;
wire [1508:0] c_w_1114;
wire [1508:0] c_w_1115;
wire [1508:0] c_w_1116;
wire [1508:0] c_w_1117;
wire [1508:0] c_w_1118;
wire [1508:0] c_w_1119;
wire [1508:0] c_w_1120;
wire [1508:0] c_w_1121;
wire [1508:0] c_w_1122;
wire [1508:0] c_w_1123;
wire [1508:0] c_w_1124;
wire [1508:0] c_w_1125;
wire [1508:0] c_w_1126;
wire [1508:0] c_w_1127;
wire [1508:0] c_w_1128;
wire [1508:0] c_w_1129;
wire [1508:0] c_w_1130;
wire [1508:0] c_w_1131;
wire [1508:0] c_w_1132;
wire [1508:0] c_w_1133;
wire [1508:0] c_w_1134;
wire [1508:0] c_w_1135;
wire [1508:0] c_w_1136;
wire [1508:0] c_w_1137;
wire [1508:0] c_w_1138;
wire [1508:0] c_w_1139;
wire [1508:0] c_w_1140;
wire [1508:0] c_w_1141;
wire [1508:0] c_w_1142;
wire [1508:0] c_w_1143;
wire [1508:0] c_w_1144;
wire [1508:0] c_w_1145;
wire [1508:0] c_w_1146;
wire [1508:0] c_w_1147;
wire [1508:0] c_w_1148;
wire [1508:0] c_w_1149;
wire [1508:0] c_w_1150;
wire [1508:0] c_w_1151;
wire [1508:0] c_w_1152;
wire [1508:0] c_w_1153;
wire [1508:0] c_w_1154;
wire [1508:0] c_w_1155;
wire [1508:0] c_w_1156;
wire [1508:0] c_w_1157;
wire [1508:0] c_w_1158;
wire [1508:0] c_w_1159;
wire [1508:0] c_w_1160;
wire [1508:0] c_w_1161;
wire [1508:0] c_w_1162;
wire [1508:0] c_w_1163;
wire [1508:0] c_w_1164;
wire [1508:0] c_w_1165;
wire [1508:0] c_w_1166;
wire [1508:0] c_w_1167;
wire [1508:0] c_w_1168;
wire [1508:0] c_w_1169;
wire [1508:0] c_w_1170;
wire [1508:0] c_w_1171;
wire [1508:0] c_w_1172;
wire [1508:0] c_w_1173;
wire [1508:0] c_w_1174;
wire [1508:0] c_w_1175;
wire [1508:0] c_w_1176;
wire [1508:0] c_w_1177;
wire [1508:0] c_w_1178;
wire [1508:0] c_w_1179;
wire [1508:0] c_w_1180;
wire [1508:0] c_w_1181;
wire [1508:0] c_w_1182;
wire [1508:0] c_w_1183;
wire [1508:0] c_w_1184;
wire [1508:0] c_w_1185;
wire [1508:0] c_w_1186;
wire [1508:0] c_w_1187;
wire [1508:0] c_w_1188;
wire [1508:0] c_w_1189;
wire [1508:0] c_w_1190;
wire [1508:0] c_w_1191;
wire [1508:0] c_w_1192;
wire [1508:0] c_w_1193;
wire [1508:0] c_w_1194;
wire [1508:0] c_w_1195;
wire [1508:0] c_w_1196;
wire [1508:0] c_w_1197;
wire [1508:0] c_w_1198;
wire [1508:0] c_w_1199;
wire [1508:0] c_w_1200;
wire [1508:0] c_w_1201;
wire [1508:0] c_w_1202;
wire [1508:0] c_w_1203;
wire [1508:0] c_w_1204;
wire [1508:0] c_w_1205;
wire [1508:0] c_w_1206;
wire [1508:0] c_w_1207;
wire [1508:0] c_w_1208;
wire [1508:0] c_w_1209;
wire [1508:0] c_w_1210;
wire [1508:0] c_w_1211;
wire [1508:0] c_w_1212;
wire [1508:0] c_w_1213;
wire [1508:0] c_w_1214;
wire [1508:0] c_w_1215;
wire [1508:0] c_w_1216;
wire [1508:0] c_w_1217;
wire [1508:0] c_w_1218;
wire [1508:0] c_w_1219;
wire [1508:0] c_w_1220;
wire [1508:0] c_w_1221;
wire [1508:0] c_w_1222;
wire [1508:0] c_w_1223;
wire [1508:0] c_w_1224;
wire [1508:0] c_w_1225;
wire [1508:0] c_w_1226;
wire [1508:0] c_w_1227;
wire [1508:0] c_w_1228;
wire [1508:0] c_w_1229;
wire [1508:0] c_w_1230;
wire [1508:0] c_w_1231;
wire [1508:0] c_w_1232;
wire [1508:0] c_w_1233;
wire [1508:0] c_w_1234;
wire [1508:0] c_w_1235;
wire [1508:0] c_w_1236;
wire [1508:0] c_w_1237;
wire [1508:0] c_w_1238;
wire [1508:0] c_w_1239;
wire [1508:0] c_w_1240;
wire [1508:0] c_w_1241;
wire [1508:0] c_w_1242;
wire [1508:0] c_w_1243;
wire [1508:0] c_w_1244;
wire [1508:0] c_w_1245;
wire [1508:0] c_w_1246;
wire [1508:0] c_w_1247;
wire [1508:0] c_w_1248;
wire [1508:0] c_w_1249;
wire [1508:0] c_w_1250;
wire [1508:0] c_w_1251;
wire [1508:0] c_w_1252;
wire [1508:0] c_w_1253;
wire [1508:0] c_w_1254;
wire [1508:0] c_w_1255;
wire [1508:0] c_w_1256;
wire [1508:0] c_w_1257;
wire [1508:0] c_w_1258;
wire [1508:0] c_w_1259;
wire [1508:0] c_w_1260;
wire [1508:0] c_w_1261;
wire [1508:0] c_w_1262;
wire [1508:0] c_w_1263;
wire [1508:0] c_w_1264;
wire [1508:0] c_w_1265;
wire [1508:0] c_w_1266;
wire [1508:0] c_w_1267;
wire [1508:0] c_w_1268;
wire [1508:0] c_w_1269;
wire [1508:0] c_w_1270;
wire [1508:0] c_w_1271;
wire [1508:0] c_w_1272;
wire [1508:0] c_w_1273;
wire [1508:0] c_w_1274;
wire [1508:0] c_w_1275;
wire [1508:0] c_w_1276;
wire [1508:0] c_w_1277;
wire [1508:0] c_w_1278;
wire [1508:0] c_w_1279;
wire [1508:0] c_w_1280;
wire [1508:0] c_w_1281;
wire [1508:0] c_w_1282;
wire [1508:0] c_w_1283;
wire [1508:0] c_w_1284;
wire [1508:0] c_w_1285;
wire [1508:0] c_w_1286;
wire [1508:0] c_w_1287;
wire [1508:0] c_w_1288;
wire [1508:0] c_w_1289;
wire [1508:0] c_w_1290;
wire [1508:0] c_w_1291;
wire [1508:0] c_w_1292;
wire [1508:0] c_w_1293;
wire [1508:0] c_w_1294;
wire [1508:0] c_w_1295;
wire [1508:0] c_w_1296;
wire [1508:0] c_w_1297;
wire [1508:0] c_w_1298;
wire [1508:0] c_w_1299;
wire [1508:0] c_w_1300;
wire [1508:0] c_w_1301;
wire [1508:0] c_w_1302;
wire [1508:0] c_w_1303;
wire [1508:0] c_w_1304;
wire [1508:0] c_w_1305;
wire [1508:0] c_w_1306;
wire [1508:0] c_w_1307;
wire [1508:0] c_w_1308;
wire [1508:0] c_w_1309;
wire [1508:0] c_w_1310;
wire [1508:0] c_w_1311;
wire [1508:0] c_w_1312;
wire [1508:0] c_w_1313;
wire [1508:0] c_w_1314;
wire [1508:0] c_w_1315;
wire [1508:0] c_w_1316;
wire [1508:0] c_w_1317;
wire [1508:0] c_w_1318;
wire [1508:0] c_w_1319;
wire [1508:0] c_w_1320;
wire [1508:0] c_w_1321;
wire [1508:0] c_w_1322;
wire [1508:0] c_w_1323;
wire [1508:0] c_w_1324;
wire [1508:0] c_w_1325;
wire [1508:0] c_w_1326;
wire [1508:0] c_w_1327;
wire [1508:0] c_w_1328;
wire [1508:0] c_w_1329;
wire [1508:0] c_w_1330;
wire [1508:0] c_w_1331;
wire [1508:0] c_w_1332;
wire [1508:0] c_w_1333;
wire [1508:0] c_w_1334;
wire [1508:0] c_w_1335;
wire [1508:0] c_w_1336;
wire [1508:0] c_w_1337;
wire [1508:0] c_w_1338;
wire [1508:0] c_w_1339;
wire [1508:0] c_w_1340;
wire [1508:0] c_w_1341;
wire [1508:0] c_w_1342;
wire [1508:0] c_w_1343;
wire [1508:0] c_w_1344;
wire [1508:0] c_w_1345;
wire [1508:0] c_w_1346;
wire [1508:0] c_w_1347;
wire [1508:0] c_w_1348;
wire [1508:0] c_w_1349;
wire [1508:0] c_w_1350;
wire [1508:0] c_w_1351;
wire [1508:0] c_w_1352;
wire [1508:0] c_w_1353;
wire [1508:0] c_w_1354;
wire [1508:0] c_w_1355;
wire [1508:0] c_w_1356;
wire [1508:0] c_w_1357;
wire [1508:0] c_w_1358;
wire [1508:0] c_w_1359;
wire [1508:0] c_w_1360;
wire [1508:0] c_w_1361;
wire [1508:0] c_w_1362;
wire [1508:0] c_w_1363;
wire [1508:0] c_w_1364;
wire [1508:0] c_w_1365;
wire [1508:0] c_w_1366;
wire [1508:0] c_w_1367;
wire [1508:0] c_w_1368;
wire [1508:0] c_w_1369;
wire [1508:0] c_w_1370;
wire [1508:0] c_w_1371;
wire [1508:0] c_w_1372;
wire [1508:0] c_w_1373;
wire [1508:0] c_w_1374;
wire [1508:0] c_w_1375;
wire [1508:0] c_w_1376;
wire [1508:0] c_w_1377;
wire [1508:0] c_w_1378;
wire [1508:0] c_w_1379;
wire [1508:0] c_w_1380;
wire [1508:0] c_w_1381;
wire [1508:0] c_w_1382;
wire [1508:0] c_w_1383;
wire [1508:0] c_w_1384;
wire [1508:0] c_w_1385;
wire [1508:0] c_w_1386;
wire [1508:0] c_w_1387;
wire [1508:0] c_w_1388;
wire [1508:0] c_w_1389;
wire [1508:0] c_w_1390;
wire [1508:0] c_w_1391;
wire [1508:0] c_w_1392;
wire [1508:0] c_w_1393;
wire [1508:0] c_w_1394;
wire [1508:0] c_w_1395;
wire [1508:0] c_w_1396;
wire [1508:0] c_w_1397;
wire [1508:0] c_w_1398;
wire [1508:0] c_w_1399;
wire [1508:0] c_w_1400;
wire [1508:0] c_w_1401;
wire [1508:0] c_w_1402;
wire [1508:0] c_w_1403;
wire [1508:0] c_w_1404;
wire [1508:0] c_w_1405;
wire [1508:0] c_w_1406;
wire [1508:0] c_w_1407;
wire [1508:0] c_w_1408;
wire [1508:0] c_w_1409;
wire [1508:0] c_w_1410;
wire [1508:0] c_w_1411;
wire [1508:0] c_w_1412;
wire [1508:0] c_w_1413;
wire [1508:0] c_w_1414;
wire [1508:0] c_w_1415;
wire [1508:0] c_w_1416;
wire [1508:0] c_w_1417;
wire [1508:0] c_w_1418;
wire [1508:0] c_w_1419;
wire [1508:0] c_w_1420;
wire [1508:0] c_w_1421;
wire [1508:0] c_w_1422;
wire [1508:0] c_w_1423;
wire [1508:0] c_w_1424;
wire [1508:0] c_w_1425;
wire [1508:0] c_w_1426;
wire [1508:0] c_w_1427;
wire [1508:0] c_w_1428;
wire [1508:0] c_w_1429;
wire [1508:0] c_w_1430;
wire [1508:0] c_w_1431;
wire [1508:0] c_w_1432;
wire [1508:0] c_w_1433;
wire [1508:0] c_w_1434;
wire [1508:0] c_w_1435;
wire [1508:0] c_w_1436;
wire [1508:0] c_w_1437;
wire [1508:0] c_w_1438;
wire [1508:0] c_w_1439;
wire [1508:0] c_w_1440;
wire [1508:0] c_w_1441;
wire [1508:0] c_w_1442;
wire [1508:0] c_w_1443;
wire [1508:0] c_w_1444;
wire [1508:0] c_w_1445;
wire [1508:0] c_w_1446;
wire [1508:0] c_w_1447;
wire [1508:0] c_w_1448;
wire [1508:0] c_w_1449;
wire [1508:0] c_w_1450;
wire [1508:0] c_w_1451;
wire [1508:0] c_w_1452;
wire [1508:0] c_w_1453;
wire [1508:0] c_w_1454;
wire [1508:0] c_w_1455;
wire [1508:0] c_w_1456;
wire [1508:0] c_w_1457;
wire [1508:0] c_w_1458;
wire [1508:0] c_w_1459;
wire [1508:0] c_w_1460;
wire [1508:0] c_w_1461;
wire [1508:0] c_w_1462;
wire [1508:0] c_w_1463;
wire [1508:0] c_w_1464;
wire [1508:0] c_w_1465;
wire [1508:0] c_w_1466;
wire [1508:0] c_w_1467;
wire [1508:0] c_w_1468;
wire [1508:0] c_w_1469;
wire [1508:0] c_w_1470;
wire [1508:0] c_w_1471;
wire [1508:0] c_w_1472;
wire [1508:0] c_w_1473;
wire [1508:0] c_w_1474;
wire [1508:0] c_w_1475;
wire [1508:0] c_w_1476;
wire [1508:0] c_w_1477;
wire [1508:0] c_w_1478;
wire [1508:0] c_w_1479;
wire [1508:0] c_w_1480;
wire [1508:0] c_w_1481;
wire [1508:0] c_w_1482;
wire [1508:0] c_w_1483;
wire [1508:0] c_w_1484;
wire [1508:0] c_w_1485;
wire [1508:0] c_w_1486;
wire [1508:0] c_w_1487;
wire [1508:0] c_w_1488;
wire [1508:0] c_w_1489;
wire [1508:0] c_w_1490;
wire [1508:0] c_w_1491;
wire [1508:0] c_w_1492;
wire [1508:0] c_w_1493;
wire [1508:0] c_w_1494;
wire [1508:0] c_w_1495;
wire [1508:0] c_w_1496;
wire [1508:0] c_w_1497;
wire [1508:0] c_w_1498;
wire [1508:0] c_w_1499;
wire [1508:0] c_w_1500;
wire [1508:0] c_w_1501;
wire [1508:0] c_w_1502;
wire [1508:0] c_w_1503;
wire [1508:0] c_w_1504;
wire [1508:0] c_w_1505;
wire [1508:0] c_w_1506;
wire [1508:0] c_w_1507;
wire [1508:0] c_w_1508;
    
AND_array_1509 AND_array_1509_i0(a,b[0],c_w_0);
AND_array_1509 AND_array_1509_i1(a,b[1],c_w_1);
AND_array_1509 AND_array_1509_i2(a,b[2],c_w_2);
AND_array_1509 AND_array_1509_i3(a,b[3],c_w_3);
AND_array_1509 AND_array_1509_i4(a,b[4],c_w_4);
AND_array_1509 AND_array_1509_i5(a,b[5],c_w_5);
AND_array_1509 AND_array_1509_i6(a,b[6],c_w_6);
AND_array_1509 AND_array_1509_i7(a,b[7],c_w_7);
AND_array_1509 AND_array_1509_i8(a,b[8],c_w_8);
AND_array_1509 AND_array_1509_i9(a,b[9],c_w_9);
AND_array_1509 AND_array_1509_i10(a,b[10],c_w_10);
AND_array_1509 AND_array_1509_i11(a,b[11],c_w_11);
AND_array_1509 AND_array_1509_i12(a,b[12],c_w_12);
AND_array_1509 AND_array_1509_i13(a,b[13],c_w_13);
AND_array_1509 AND_array_1509_i14(a,b[14],c_w_14);
AND_array_1509 AND_array_1509_i15(a,b[15],c_w_15);
AND_array_1509 AND_array_1509_i16(a,b[16],c_w_16);
AND_array_1509 AND_array_1509_i17(a,b[17],c_w_17);
AND_array_1509 AND_array_1509_i18(a,b[18],c_w_18);
AND_array_1509 AND_array_1509_i19(a,b[19],c_w_19);
AND_array_1509 AND_array_1509_i20(a,b[20],c_w_20);
AND_array_1509 AND_array_1509_i21(a,b[21],c_w_21);
AND_array_1509 AND_array_1509_i22(a,b[22],c_w_22);
AND_array_1509 AND_array_1509_i23(a,b[23],c_w_23);
AND_array_1509 AND_array_1509_i24(a,b[24],c_w_24);
AND_array_1509 AND_array_1509_i25(a,b[25],c_w_25);
AND_array_1509 AND_array_1509_i26(a,b[26],c_w_26);
AND_array_1509 AND_array_1509_i27(a,b[27],c_w_27);
AND_array_1509 AND_array_1509_i28(a,b[28],c_w_28);
AND_array_1509 AND_array_1509_i29(a,b[29],c_w_29);
AND_array_1509 AND_array_1509_i30(a,b[30],c_w_30);
AND_array_1509 AND_array_1509_i31(a,b[31],c_w_31);
AND_array_1509 AND_array_1509_i32(a,b[32],c_w_32);
AND_array_1509 AND_array_1509_i33(a,b[33],c_w_33);
AND_array_1509 AND_array_1509_i34(a,b[34],c_w_34);
AND_array_1509 AND_array_1509_i35(a,b[35],c_w_35);
AND_array_1509 AND_array_1509_i36(a,b[36],c_w_36);
AND_array_1509 AND_array_1509_i37(a,b[37],c_w_37);
AND_array_1509 AND_array_1509_i38(a,b[38],c_w_38);
AND_array_1509 AND_array_1509_i39(a,b[39],c_w_39);
AND_array_1509 AND_array_1509_i40(a,b[40],c_w_40);
AND_array_1509 AND_array_1509_i41(a,b[41],c_w_41);
AND_array_1509 AND_array_1509_i42(a,b[42],c_w_42);
AND_array_1509 AND_array_1509_i43(a,b[43],c_w_43);
AND_array_1509 AND_array_1509_i44(a,b[44],c_w_44);
AND_array_1509 AND_array_1509_i45(a,b[45],c_w_45);
AND_array_1509 AND_array_1509_i46(a,b[46],c_w_46);
AND_array_1509 AND_array_1509_i47(a,b[47],c_w_47);
AND_array_1509 AND_array_1509_i48(a,b[48],c_w_48);
AND_array_1509 AND_array_1509_i49(a,b[49],c_w_49);
AND_array_1509 AND_array_1509_i50(a,b[50],c_w_50);
AND_array_1509 AND_array_1509_i51(a,b[51],c_w_51);
AND_array_1509 AND_array_1509_i52(a,b[52],c_w_52);
AND_array_1509 AND_array_1509_i53(a,b[53],c_w_53);
AND_array_1509 AND_array_1509_i54(a,b[54],c_w_54);
AND_array_1509 AND_array_1509_i55(a,b[55],c_w_55);
AND_array_1509 AND_array_1509_i56(a,b[56],c_w_56);
AND_array_1509 AND_array_1509_i57(a,b[57],c_w_57);
AND_array_1509 AND_array_1509_i58(a,b[58],c_w_58);
AND_array_1509 AND_array_1509_i59(a,b[59],c_w_59);
AND_array_1509 AND_array_1509_i60(a,b[60],c_w_60);
AND_array_1509 AND_array_1509_i61(a,b[61],c_w_61);
AND_array_1509 AND_array_1509_i62(a,b[62],c_w_62);
AND_array_1509 AND_array_1509_i63(a,b[63],c_w_63);
AND_array_1509 AND_array_1509_i64(a,b[64],c_w_64);
AND_array_1509 AND_array_1509_i65(a,b[65],c_w_65);
AND_array_1509 AND_array_1509_i66(a,b[66],c_w_66);
AND_array_1509 AND_array_1509_i67(a,b[67],c_w_67);
AND_array_1509 AND_array_1509_i68(a,b[68],c_w_68);
AND_array_1509 AND_array_1509_i69(a,b[69],c_w_69);
AND_array_1509 AND_array_1509_i70(a,b[70],c_w_70);
AND_array_1509 AND_array_1509_i71(a,b[71],c_w_71);
AND_array_1509 AND_array_1509_i72(a,b[72],c_w_72);
AND_array_1509 AND_array_1509_i73(a,b[73],c_w_73);
AND_array_1509 AND_array_1509_i74(a,b[74],c_w_74);
AND_array_1509 AND_array_1509_i75(a,b[75],c_w_75);
AND_array_1509 AND_array_1509_i76(a,b[76],c_w_76);
AND_array_1509 AND_array_1509_i77(a,b[77],c_w_77);
AND_array_1509 AND_array_1509_i78(a,b[78],c_w_78);
AND_array_1509 AND_array_1509_i79(a,b[79],c_w_79);
AND_array_1509 AND_array_1509_i80(a,b[80],c_w_80);
AND_array_1509 AND_array_1509_i81(a,b[81],c_w_81);
AND_array_1509 AND_array_1509_i82(a,b[82],c_w_82);
AND_array_1509 AND_array_1509_i83(a,b[83],c_w_83);
AND_array_1509 AND_array_1509_i84(a,b[84],c_w_84);
AND_array_1509 AND_array_1509_i85(a,b[85],c_w_85);
AND_array_1509 AND_array_1509_i86(a,b[86],c_w_86);
AND_array_1509 AND_array_1509_i87(a,b[87],c_w_87);
AND_array_1509 AND_array_1509_i88(a,b[88],c_w_88);
AND_array_1509 AND_array_1509_i89(a,b[89],c_w_89);
AND_array_1509 AND_array_1509_i90(a,b[90],c_w_90);
AND_array_1509 AND_array_1509_i91(a,b[91],c_w_91);
AND_array_1509 AND_array_1509_i92(a,b[92],c_w_92);
AND_array_1509 AND_array_1509_i93(a,b[93],c_w_93);
AND_array_1509 AND_array_1509_i94(a,b[94],c_w_94);
AND_array_1509 AND_array_1509_i95(a,b[95],c_w_95);
AND_array_1509 AND_array_1509_i96(a,b[96],c_w_96);
AND_array_1509 AND_array_1509_i97(a,b[97],c_w_97);
AND_array_1509 AND_array_1509_i98(a,b[98],c_w_98);
AND_array_1509 AND_array_1509_i99(a,b[99],c_w_99);
AND_array_1509 AND_array_1509_i100(a,b[100],c_w_100);
AND_array_1509 AND_array_1509_i101(a,b[101],c_w_101);
AND_array_1509 AND_array_1509_i102(a,b[102],c_w_102);
AND_array_1509 AND_array_1509_i103(a,b[103],c_w_103);
AND_array_1509 AND_array_1509_i104(a,b[104],c_w_104);
AND_array_1509 AND_array_1509_i105(a,b[105],c_w_105);
AND_array_1509 AND_array_1509_i106(a,b[106],c_w_106);
AND_array_1509 AND_array_1509_i107(a,b[107],c_w_107);
AND_array_1509 AND_array_1509_i108(a,b[108],c_w_108);
AND_array_1509 AND_array_1509_i109(a,b[109],c_w_109);
AND_array_1509 AND_array_1509_i110(a,b[110],c_w_110);
AND_array_1509 AND_array_1509_i111(a,b[111],c_w_111);
AND_array_1509 AND_array_1509_i112(a,b[112],c_w_112);
AND_array_1509 AND_array_1509_i113(a,b[113],c_w_113);
AND_array_1509 AND_array_1509_i114(a,b[114],c_w_114);
AND_array_1509 AND_array_1509_i115(a,b[115],c_w_115);
AND_array_1509 AND_array_1509_i116(a,b[116],c_w_116);
AND_array_1509 AND_array_1509_i117(a,b[117],c_w_117);
AND_array_1509 AND_array_1509_i118(a,b[118],c_w_118);
AND_array_1509 AND_array_1509_i119(a,b[119],c_w_119);
AND_array_1509 AND_array_1509_i120(a,b[120],c_w_120);
AND_array_1509 AND_array_1509_i121(a,b[121],c_w_121);
AND_array_1509 AND_array_1509_i122(a,b[122],c_w_122);
AND_array_1509 AND_array_1509_i123(a,b[123],c_w_123);
AND_array_1509 AND_array_1509_i124(a,b[124],c_w_124);
AND_array_1509 AND_array_1509_i125(a,b[125],c_w_125);
AND_array_1509 AND_array_1509_i126(a,b[126],c_w_126);
AND_array_1509 AND_array_1509_i127(a,b[127],c_w_127);
AND_array_1509 AND_array_1509_i128(a,b[128],c_w_128);
AND_array_1509 AND_array_1509_i129(a,b[129],c_w_129);
AND_array_1509 AND_array_1509_i130(a,b[130],c_w_130);
AND_array_1509 AND_array_1509_i131(a,b[131],c_w_131);
AND_array_1509 AND_array_1509_i132(a,b[132],c_w_132);
AND_array_1509 AND_array_1509_i133(a,b[133],c_w_133);
AND_array_1509 AND_array_1509_i134(a,b[134],c_w_134);
AND_array_1509 AND_array_1509_i135(a,b[135],c_w_135);
AND_array_1509 AND_array_1509_i136(a,b[136],c_w_136);
AND_array_1509 AND_array_1509_i137(a,b[137],c_w_137);
AND_array_1509 AND_array_1509_i138(a,b[138],c_w_138);
AND_array_1509 AND_array_1509_i139(a,b[139],c_w_139);
AND_array_1509 AND_array_1509_i140(a,b[140],c_w_140);
AND_array_1509 AND_array_1509_i141(a,b[141],c_w_141);
AND_array_1509 AND_array_1509_i142(a,b[142],c_w_142);
AND_array_1509 AND_array_1509_i143(a,b[143],c_w_143);
AND_array_1509 AND_array_1509_i144(a,b[144],c_w_144);
AND_array_1509 AND_array_1509_i145(a,b[145],c_w_145);
AND_array_1509 AND_array_1509_i146(a,b[146],c_w_146);
AND_array_1509 AND_array_1509_i147(a,b[147],c_w_147);
AND_array_1509 AND_array_1509_i148(a,b[148],c_w_148);
AND_array_1509 AND_array_1509_i149(a,b[149],c_w_149);
AND_array_1509 AND_array_1509_i150(a,b[150],c_w_150);
AND_array_1509 AND_array_1509_i151(a,b[151],c_w_151);
AND_array_1509 AND_array_1509_i152(a,b[152],c_w_152);
AND_array_1509 AND_array_1509_i153(a,b[153],c_w_153);
AND_array_1509 AND_array_1509_i154(a,b[154],c_w_154);
AND_array_1509 AND_array_1509_i155(a,b[155],c_w_155);
AND_array_1509 AND_array_1509_i156(a,b[156],c_w_156);
AND_array_1509 AND_array_1509_i157(a,b[157],c_w_157);
AND_array_1509 AND_array_1509_i158(a,b[158],c_w_158);
AND_array_1509 AND_array_1509_i159(a,b[159],c_w_159);
AND_array_1509 AND_array_1509_i160(a,b[160],c_w_160);
AND_array_1509 AND_array_1509_i161(a,b[161],c_w_161);
AND_array_1509 AND_array_1509_i162(a,b[162],c_w_162);
AND_array_1509 AND_array_1509_i163(a,b[163],c_w_163);
AND_array_1509 AND_array_1509_i164(a,b[164],c_w_164);
AND_array_1509 AND_array_1509_i165(a,b[165],c_w_165);
AND_array_1509 AND_array_1509_i166(a,b[166],c_w_166);
AND_array_1509 AND_array_1509_i167(a,b[167],c_w_167);
AND_array_1509 AND_array_1509_i168(a,b[168],c_w_168);
AND_array_1509 AND_array_1509_i169(a,b[169],c_w_169);
AND_array_1509 AND_array_1509_i170(a,b[170],c_w_170);
AND_array_1509 AND_array_1509_i171(a,b[171],c_w_171);
AND_array_1509 AND_array_1509_i172(a,b[172],c_w_172);
AND_array_1509 AND_array_1509_i173(a,b[173],c_w_173);
AND_array_1509 AND_array_1509_i174(a,b[174],c_w_174);
AND_array_1509 AND_array_1509_i175(a,b[175],c_w_175);
AND_array_1509 AND_array_1509_i176(a,b[176],c_w_176);
AND_array_1509 AND_array_1509_i177(a,b[177],c_w_177);
AND_array_1509 AND_array_1509_i178(a,b[178],c_w_178);
AND_array_1509 AND_array_1509_i179(a,b[179],c_w_179);
AND_array_1509 AND_array_1509_i180(a,b[180],c_w_180);
AND_array_1509 AND_array_1509_i181(a,b[181],c_w_181);
AND_array_1509 AND_array_1509_i182(a,b[182],c_w_182);
AND_array_1509 AND_array_1509_i183(a,b[183],c_w_183);
AND_array_1509 AND_array_1509_i184(a,b[184],c_w_184);
AND_array_1509 AND_array_1509_i185(a,b[185],c_w_185);
AND_array_1509 AND_array_1509_i186(a,b[186],c_w_186);
AND_array_1509 AND_array_1509_i187(a,b[187],c_w_187);
AND_array_1509 AND_array_1509_i188(a,b[188],c_w_188);
AND_array_1509 AND_array_1509_i189(a,b[189],c_w_189);
AND_array_1509 AND_array_1509_i190(a,b[190],c_w_190);
AND_array_1509 AND_array_1509_i191(a,b[191],c_w_191);
AND_array_1509 AND_array_1509_i192(a,b[192],c_w_192);
AND_array_1509 AND_array_1509_i193(a,b[193],c_w_193);
AND_array_1509 AND_array_1509_i194(a,b[194],c_w_194);
AND_array_1509 AND_array_1509_i195(a,b[195],c_w_195);
AND_array_1509 AND_array_1509_i196(a,b[196],c_w_196);
AND_array_1509 AND_array_1509_i197(a,b[197],c_w_197);
AND_array_1509 AND_array_1509_i198(a,b[198],c_w_198);
AND_array_1509 AND_array_1509_i199(a,b[199],c_w_199);
AND_array_1509 AND_array_1509_i200(a,b[200],c_w_200);
AND_array_1509 AND_array_1509_i201(a,b[201],c_w_201);
AND_array_1509 AND_array_1509_i202(a,b[202],c_w_202);
AND_array_1509 AND_array_1509_i203(a,b[203],c_w_203);
AND_array_1509 AND_array_1509_i204(a,b[204],c_w_204);
AND_array_1509 AND_array_1509_i205(a,b[205],c_w_205);
AND_array_1509 AND_array_1509_i206(a,b[206],c_w_206);
AND_array_1509 AND_array_1509_i207(a,b[207],c_w_207);
AND_array_1509 AND_array_1509_i208(a,b[208],c_w_208);
AND_array_1509 AND_array_1509_i209(a,b[209],c_w_209);
AND_array_1509 AND_array_1509_i210(a,b[210],c_w_210);
AND_array_1509 AND_array_1509_i211(a,b[211],c_w_211);
AND_array_1509 AND_array_1509_i212(a,b[212],c_w_212);
AND_array_1509 AND_array_1509_i213(a,b[213],c_w_213);
AND_array_1509 AND_array_1509_i214(a,b[214],c_w_214);
AND_array_1509 AND_array_1509_i215(a,b[215],c_w_215);
AND_array_1509 AND_array_1509_i216(a,b[216],c_w_216);
AND_array_1509 AND_array_1509_i217(a,b[217],c_w_217);
AND_array_1509 AND_array_1509_i218(a,b[218],c_w_218);
AND_array_1509 AND_array_1509_i219(a,b[219],c_w_219);
AND_array_1509 AND_array_1509_i220(a,b[220],c_w_220);
AND_array_1509 AND_array_1509_i221(a,b[221],c_w_221);
AND_array_1509 AND_array_1509_i222(a,b[222],c_w_222);
AND_array_1509 AND_array_1509_i223(a,b[223],c_w_223);
AND_array_1509 AND_array_1509_i224(a,b[224],c_w_224);
AND_array_1509 AND_array_1509_i225(a,b[225],c_w_225);
AND_array_1509 AND_array_1509_i226(a,b[226],c_w_226);
AND_array_1509 AND_array_1509_i227(a,b[227],c_w_227);
AND_array_1509 AND_array_1509_i228(a,b[228],c_w_228);
AND_array_1509 AND_array_1509_i229(a,b[229],c_w_229);
AND_array_1509 AND_array_1509_i230(a,b[230],c_w_230);
AND_array_1509 AND_array_1509_i231(a,b[231],c_w_231);
AND_array_1509 AND_array_1509_i232(a,b[232],c_w_232);
AND_array_1509 AND_array_1509_i233(a,b[233],c_w_233);
AND_array_1509 AND_array_1509_i234(a,b[234],c_w_234);
AND_array_1509 AND_array_1509_i235(a,b[235],c_w_235);
AND_array_1509 AND_array_1509_i236(a,b[236],c_w_236);
AND_array_1509 AND_array_1509_i237(a,b[237],c_w_237);
AND_array_1509 AND_array_1509_i238(a,b[238],c_w_238);
AND_array_1509 AND_array_1509_i239(a,b[239],c_w_239);
AND_array_1509 AND_array_1509_i240(a,b[240],c_w_240);
AND_array_1509 AND_array_1509_i241(a,b[241],c_w_241);
AND_array_1509 AND_array_1509_i242(a,b[242],c_w_242);
AND_array_1509 AND_array_1509_i243(a,b[243],c_w_243);
AND_array_1509 AND_array_1509_i244(a,b[244],c_w_244);
AND_array_1509 AND_array_1509_i245(a,b[245],c_w_245);
AND_array_1509 AND_array_1509_i246(a,b[246],c_w_246);
AND_array_1509 AND_array_1509_i247(a,b[247],c_w_247);
AND_array_1509 AND_array_1509_i248(a,b[248],c_w_248);
AND_array_1509 AND_array_1509_i249(a,b[249],c_w_249);
AND_array_1509 AND_array_1509_i250(a,b[250],c_w_250);
AND_array_1509 AND_array_1509_i251(a,b[251],c_w_251);
AND_array_1509 AND_array_1509_i252(a,b[252],c_w_252);
AND_array_1509 AND_array_1509_i253(a,b[253],c_w_253);
AND_array_1509 AND_array_1509_i254(a,b[254],c_w_254);
AND_array_1509 AND_array_1509_i255(a,b[255],c_w_255);
AND_array_1509 AND_array_1509_i256(a,b[256],c_w_256);
AND_array_1509 AND_array_1509_i257(a,b[257],c_w_257);
AND_array_1509 AND_array_1509_i258(a,b[258],c_w_258);
AND_array_1509 AND_array_1509_i259(a,b[259],c_w_259);
AND_array_1509 AND_array_1509_i260(a,b[260],c_w_260);
AND_array_1509 AND_array_1509_i261(a,b[261],c_w_261);
AND_array_1509 AND_array_1509_i262(a,b[262],c_w_262);
AND_array_1509 AND_array_1509_i263(a,b[263],c_w_263);
AND_array_1509 AND_array_1509_i264(a,b[264],c_w_264);
AND_array_1509 AND_array_1509_i265(a,b[265],c_w_265);
AND_array_1509 AND_array_1509_i266(a,b[266],c_w_266);
AND_array_1509 AND_array_1509_i267(a,b[267],c_w_267);
AND_array_1509 AND_array_1509_i268(a,b[268],c_w_268);
AND_array_1509 AND_array_1509_i269(a,b[269],c_w_269);
AND_array_1509 AND_array_1509_i270(a,b[270],c_w_270);
AND_array_1509 AND_array_1509_i271(a,b[271],c_w_271);
AND_array_1509 AND_array_1509_i272(a,b[272],c_w_272);
AND_array_1509 AND_array_1509_i273(a,b[273],c_w_273);
AND_array_1509 AND_array_1509_i274(a,b[274],c_w_274);
AND_array_1509 AND_array_1509_i275(a,b[275],c_w_275);
AND_array_1509 AND_array_1509_i276(a,b[276],c_w_276);
AND_array_1509 AND_array_1509_i277(a,b[277],c_w_277);
AND_array_1509 AND_array_1509_i278(a,b[278],c_w_278);
AND_array_1509 AND_array_1509_i279(a,b[279],c_w_279);
AND_array_1509 AND_array_1509_i280(a,b[280],c_w_280);
AND_array_1509 AND_array_1509_i281(a,b[281],c_w_281);
AND_array_1509 AND_array_1509_i282(a,b[282],c_w_282);
AND_array_1509 AND_array_1509_i283(a,b[283],c_w_283);
AND_array_1509 AND_array_1509_i284(a,b[284],c_w_284);
AND_array_1509 AND_array_1509_i285(a,b[285],c_w_285);
AND_array_1509 AND_array_1509_i286(a,b[286],c_w_286);
AND_array_1509 AND_array_1509_i287(a,b[287],c_w_287);
AND_array_1509 AND_array_1509_i288(a,b[288],c_w_288);
AND_array_1509 AND_array_1509_i289(a,b[289],c_w_289);
AND_array_1509 AND_array_1509_i290(a,b[290],c_w_290);
AND_array_1509 AND_array_1509_i291(a,b[291],c_w_291);
AND_array_1509 AND_array_1509_i292(a,b[292],c_w_292);
AND_array_1509 AND_array_1509_i293(a,b[293],c_w_293);
AND_array_1509 AND_array_1509_i294(a,b[294],c_w_294);
AND_array_1509 AND_array_1509_i295(a,b[295],c_w_295);
AND_array_1509 AND_array_1509_i296(a,b[296],c_w_296);
AND_array_1509 AND_array_1509_i297(a,b[297],c_w_297);
AND_array_1509 AND_array_1509_i298(a,b[298],c_w_298);
AND_array_1509 AND_array_1509_i299(a,b[299],c_w_299);
AND_array_1509 AND_array_1509_i300(a,b[300],c_w_300);
AND_array_1509 AND_array_1509_i301(a,b[301],c_w_301);
AND_array_1509 AND_array_1509_i302(a,b[302],c_w_302);
AND_array_1509 AND_array_1509_i303(a,b[303],c_w_303);
AND_array_1509 AND_array_1509_i304(a,b[304],c_w_304);
AND_array_1509 AND_array_1509_i305(a,b[305],c_w_305);
AND_array_1509 AND_array_1509_i306(a,b[306],c_w_306);
AND_array_1509 AND_array_1509_i307(a,b[307],c_w_307);
AND_array_1509 AND_array_1509_i308(a,b[308],c_w_308);
AND_array_1509 AND_array_1509_i309(a,b[309],c_w_309);
AND_array_1509 AND_array_1509_i310(a,b[310],c_w_310);
AND_array_1509 AND_array_1509_i311(a,b[311],c_w_311);
AND_array_1509 AND_array_1509_i312(a,b[312],c_w_312);
AND_array_1509 AND_array_1509_i313(a,b[313],c_w_313);
AND_array_1509 AND_array_1509_i314(a,b[314],c_w_314);
AND_array_1509 AND_array_1509_i315(a,b[315],c_w_315);
AND_array_1509 AND_array_1509_i316(a,b[316],c_w_316);
AND_array_1509 AND_array_1509_i317(a,b[317],c_w_317);
AND_array_1509 AND_array_1509_i318(a,b[318],c_w_318);
AND_array_1509 AND_array_1509_i319(a,b[319],c_w_319);
AND_array_1509 AND_array_1509_i320(a,b[320],c_w_320);
AND_array_1509 AND_array_1509_i321(a,b[321],c_w_321);
AND_array_1509 AND_array_1509_i322(a,b[322],c_w_322);
AND_array_1509 AND_array_1509_i323(a,b[323],c_w_323);
AND_array_1509 AND_array_1509_i324(a,b[324],c_w_324);
AND_array_1509 AND_array_1509_i325(a,b[325],c_w_325);
AND_array_1509 AND_array_1509_i326(a,b[326],c_w_326);
AND_array_1509 AND_array_1509_i327(a,b[327],c_w_327);
AND_array_1509 AND_array_1509_i328(a,b[328],c_w_328);
AND_array_1509 AND_array_1509_i329(a,b[329],c_w_329);
AND_array_1509 AND_array_1509_i330(a,b[330],c_w_330);
AND_array_1509 AND_array_1509_i331(a,b[331],c_w_331);
AND_array_1509 AND_array_1509_i332(a,b[332],c_w_332);
AND_array_1509 AND_array_1509_i333(a,b[333],c_w_333);
AND_array_1509 AND_array_1509_i334(a,b[334],c_w_334);
AND_array_1509 AND_array_1509_i335(a,b[335],c_w_335);
AND_array_1509 AND_array_1509_i336(a,b[336],c_w_336);
AND_array_1509 AND_array_1509_i337(a,b[337],c_w_337);
AND_array_1509 AND_array_1509_i338(a,b[338],c_w_338);
AND_array_1509 AND_array_1509_i339(a,b[339],c_w_339);
AND_array_1509 AND_array_1509_i340(a,b[340],c_w_340);
AND_array_1509 AND_array_1509_i341(a,b[341],c_w_341);
AND_array_1509 AND_array_1509_i342(a,b[342],c_w_342);
AND_array_1509 AND_array_1509_i343(a,b[343],c_w_343);
AND_array_1509 AND_array_1509_i344(a,b[344],c_w_344);
AND_array_1509 AND_array_1509_i345(a,b[345],c_w_345);
AND_array_1509 AND_array_1509_i346(a,b[346],c_w_346);
AND_array_1509 AND_array_1509_i347(a,b[347],c_w_347);
AND_array_1509 AND_array_1509_i348(a,b[348],c_w_348);
AND_array_1509 AND_array_1509_i349(a,b[349],c_w_349);
AND_array_1509 AND_array_1509_i350(a,b[350],c_w_350);
AND_array_1509 AND_array_1509_i351(a,b[351],c_w_351);
AND_array_1509 AND_array_1509_i352(a,b[352],c_w_352);
AND_array_1509 AND_array_1509_i353(a,b[353],c_w_353);
AND_array_1509 AND_array_1509_i354(a,b[354],c_w_354);
AND_array_1509 AND_array_1509_i355(a,b[355],c_w_355);
AND_array_1509 AND_array_1509_i356(a,b[356],c_w_356);
AND_array_1509 AND_array_1509_i357(a,b[357],c_w_357);
AND_array_1509 AND_array_1509_i358(a,b[358],c_w_358);
AND_array_1509 AND_array_1509_i359(a,b[359],c_w_359);
AND_array_1509 AND_array_1509_i360(a,b[360],c_w_360);
AND_array_1509 AND_array_1509_i361(a,b[361],c_w_361);
AND_array_1509 AND_array_1509_i362(a,b[362],c_w_362);
AND_array_1509 AND_array_1509_i363(a,b[363],c_w_363);
AND_array_1509 AND_array_1509_i364(a,b[364],c_w_364);
AND_array_1509 AND_array_1509_i365(a,b[365],c_w_365);
AND_array_1509 AND_array_1509_i366(a,b[366],c_w_366);
AND_array_1509 AND_array_1509_i367(a,b[367],c_w_367);
AND_array_1509 AND_array_1509_i368(a,b[368],c_w_368);
AND_array_1509 AND_array_1509_i369(a,b[369],c_w_369);
AND_array_1509 AND_array_1509_i370(a,b[370],c_w_370);
AND_array_1509 AND_array_1509_i371(a,b[371],c_w_371);
AND_array_1509 AND_array_1509_i372(a,b[372],c_w_372);
AND_array_1509 AND_array_1509_i373(a,b[373],c_w_373);
AND_array_1509 AND_array_1509_i374(a,b[374],c_w_374);
AND_array_1509 AND_array_1509_i375(a,b[375],c_w_375);
AND_array_1509 AND_array_1509_i376(a,b[376],c_w_376);
AND_array_1509 AND_array_1509_i377(a,b[377],c_w_377);
AND_array_1509 AND_array_1509_i378(a,b[378],c_w_378);
AND_array_1509 AND_array_1509_i379(a,b[379],c_w_379);
AND_array_1509 AND_array_1509_i380(a,b[380],c_w_380);
AND_array_1509 AND_array_1509_i381(a,b[381],c_w_381);
AND_array_1509 AND_array_1509_i382(a,b[382],c_w_382);
AND_array_1509 AND_array_1509_i383(a,b[383],c_w_383);
AND_array_1509 AND_array_1509_i384(a,b[384],c_w_384);
AND_array_1509 AND_array_1509_i385(a,b[385],c_w_385);
AND_array_1509 AND_array_1509_i386(a,b[386],c_w_386);
AND_array_1509 AND_array_1509_i387(a,b[387],c_w_387);
AND_array_1509 AND_array_1509_i388(a,b[388],c_w_388);
AND_array_1509 AND_array_1509_i389(a,b[389],c_w_389);
AND_array_1509 AND_array_1509_i390(a,b[390],c_w_390);
AND_array_1509 AND_array_1509_i391(a,b[391],c_w_391);
AND_array_1509 AND_array_1509_i392(a,b[392],c_w_392);
AND_array_1509 AND_array_1509_i393(a,b[393],c_w_393);
AND_array_1509 AND_array_1509_i394(a,b[394],c_w_394);
AND_array_1509 AND_array_1509_i395(a,b[395],c_w_395);
AND_array_1509 AND_array_1509_i396(a,b[396],c_w_396);
AND_array_1509 AND_array_1509_i397(a,b[397],c_w_397);
AND_array_1509 AND_array_1509_i398(a,b[398],c_w_398);
AND_array_1509 AND_array_1509_i399(a,b[399],c_w_399);
AND_array_1509 AND_array_1509_i400(a,b[400],c_w_400);
AND_array_1509 AND_array_1509_i401(a,b[401],c_w_401);
AND_array_1509 AND_array_1509_i402(a,b[402],c_w_402);
AND_array_1509 AND_array_1509_i403(a,b[403],c_w_403);
AND_array_1509 AND_array_1509_i404(a,b[404],c_w_404);
AND_array_1509 AND_array_1509_i405(a,b[405],c_w_405);
AND_array_1509 AND_array_1509_i406(a,b[406],c_w_406);
AND_array_1509 AND_array_1509_i407(a,b[407],c_w_407);
AND_array_1509 AND_array_1509_i408(a,b[408],c_w_408);
AND_array_1509 AND_array_1509_i409(a,b[409],c_w_409);
AND_array_1509 AND_array_1509_i410(a,b[410],c_w_410);
AND_array_1509 AND_array_1509_i411(a,b[411],c_w_411);
AND_array_1509 AND_array_1509_i412(a,b[412],c_w_412);
AND_array_1509 AND_array_1509_i413(a,b[413],c_w_413);
AND_array_1509 AND_array_1509_i414(a,b[414],c_w_414);
AND_array_1509 AND_array_1509_i415(a,b[415],c_w_415);
AND_array_1509 AND_array_1509_i416(a,b[416],c_w_416);
AND_array_1509 AND_array_1509_i417(a,b[417],c_w_417);
AND_array_1509 AND_array_1509_i418(a,b[418],c_w_418);
AND_array_1509 AND_array_1509_i419(a,b[419],c_w_419);
AND_array_1509 AND_array_1509_i420(a,b[420],c_w_420);
AND_array_1509 AND_array_1509_i421(a,b[421],c_w_421);
AND_array_1509 AND_array_1509_i422(a,b[422],c_w_422);
AND_array_1509 AND_array_1509_i423(a,b[423],c_w_423);
AND_array_1509 AND_array_1509_i424(a,b[424],c_w_424);
AND_array_1509 AND_array_1509_i425(a,b[425],c_w_425);
AND_array_1509 AND_array_1509_i426(a,b[426],c_w_426);
AND_array_1509 AND_array_1509_i427(a,b[427],c_w_427);
AND_array_1509 AND_array_1509_i428(a,b[428],c_w_428);
AND_array_1509 AND_array_1509_i429(a,b[429],c_w_429);
AND_array_1509 AND_array_1509_i430(a,b[430],c_w_430);
AND_array_1509 AND_array_1509_i431(a,b[431],c_w_431);
AND_array_1509 AND_array_1509_i432(a,b[432],c_w_432);
AND_array_1509 AND_array_1509_i433(a,b[433],c_w_433);
AND_array_1509 AND_array_1509_i434(a,b[434],c_w_434);
AND_array_1509 AND_array_1509_i435(a,b[435],c_w_435);
AND_array_1509 AND_array_1509_i436(a,b[436],c_w_436);
AND_array_1509 AND_array_1509_i437(a,b[437],c_w_437);
AND_array_1509 AND_array_1509_i438(a,b[438],c_w_438);
AND_array_1509 AND_array_1509_i439(a,b[439],c_w_439);
AND_array_1509 AND_array_1509_i440(a,b[440],c_w_440);
AND_array_1509 AND_array_1509_i441(a,b[441],c_w_441);
AND_array_1509 AND_array_1509_i442(a,b[442],c_w_442);
AND_array_1509 AND_array_1509_i443(a,b[443],c_w_443);
AND_array_1509 AND_array_1509_i444(a,b[444],c_w_444);
AND_array_1509 AND_array_1509_i445(a,b[445],c_w_445);
AND_array_1509 AND_array_1509_i446(a,b[446],c_w_446);
AND_array_1509 AND_array_1509_i447(a,b[447],c_w_447);
AND_array_1509 AND_array_1509_i448(a,b[448],c_w_448);
AND_array_1509 AND_array_1509_i449(a,b[449],c_w_449);
AND_array_1509 AND_array_1509_i450(a,b[450],c_w_450);
AND_array_1509 AND_array_1509_i451(a,b[451],c_w_451);
AND_array_1509 AND_array_1509_i452(a,b[452],c_w_452);
AND_array_1509 AND_array_1509_i453(a,b[453],c_w_453);
AND_array_1509 AND_array_1509_i454(a,b[454],c_w_454);
AND_array_1509 AND_array_1509_i455(a,b[455],c_w_455);
AND_array_1509 AND_array_1509_i456(a,b[456],c_w_456);
AND_array_1509 AND_array_1509_i457(a,b[457],c_w_457);
AND_array_1509 AND_array_1509_i458(a,b[458],c_w_458);
AND_array_1509 AND_array_1509_i459(a,b[459],c_w_459);
AND_array_1509 AND_array_1509_i460(a,b[460],c_w_460);
AND_array_1509 AND_array_1509_i461(a,b[461],c_w_461);
AND_array_1509 AND_array_1509_i462(a,b[462],c_w_462);
AND_array_1509 AND_array_1509_i463(a,b[463],c_w_463);
AND_array_1509 AND_array_1509_i464(a,b[464],c_w_464);
AND_array_1509 AND_array_1509_i465(a,b[465],c_w_465);
AND_array_1509 AND_array_1509_i466(a,b[466],c_w_466);
AND_array_1509 AND_array_1509_i467(a,b[467],c_w_467);
AND_array_1509 AND_array_1509_i468(a,b[468],c_w_468);
AND_array_1509 AND_array_1509_i469(a,b[469],c_w_469);
AND_array_1509 AND_array_1509_i470(a,b[470],c_w_470);
AND_array_1509 AND_array_1509_i471(a,b[471],c_w_471);
AND_array_1509 AND_array_1509_i472(a,b[472],c_w_472);
AND_array_1509 AND_array_1509_i473(a,b[473],c_w_473);
AND_array_1509 AND_array_1509_i474(a,b[474],c_w_474);
AND_array_1509 AND_array_1509_i475(a,b[475],c_w_475);
AND_array_1509 AND_array_1509_i476(a,b[476],c_w_476);
AND_array_1509 AND_array_1509_i477(a,b[477],c_w_477);
AND_array_1509 AND_array_1509_i478(a,b[478],c_w_478);
AND_array_1509 AND_array_1509_i479(a,b[479],c_w_479);
AND_array_1509 AND_array_1509_i480(a,b[480],c_w_480);
AND_array_1509 AND_array_1509_i481(a,b[481],c_w_481);
AND_array_1509 AND_array_1509_i482(a,b[482],c_w_482);
AND_array_1509 AND_array_1509_i483(a,b[483],c_w_483);
AND_array_1509 AND_array_1509_i484(a,b[484],c_w_484);
AND_array_1509 AND_array_1509_i485(a,b[485],c_w_485);
AND_array_1509 AND_array_1509_i486(a,b[486],c_w_486);
AND_array_1509 AND_array_1509_i487(a,b[487],c_w_487);
AND_array_1509 AND_array_1509_i488(a,b[488],c_w_488);
AND_array_1509 AND_array_1509_i489(a,b[489],c_w_489);
AND_array_1509 AND_array_1509_i490(a,b[490],c_w_490);
AND_array_1509 AND_array_1509_i491(a,b[491],c_w_491);
AND_array_1509 AND_array_1509_i492(a,b[492],c_w_492);
AND_array_1509 AND_array_1509_i493(a,b[493],c_w_493);
AND_array_1509 AND_array_1509_i494(a,b[494],c_w_494);
AND_array_1509 AND_array_1509_i495(a,b[495],c_w_495);
AND_array_1509 AND_array_1509_i496(a,b[496],c_w_496);
AND_array_1509 AND_array_1509_i497(a,b[497],c_w_497);
AND_array_1509 AND_array_1509_i498(a,b[498],c_w_498);
AND_array_1509 AND_array_1509_i499(a,b[499],c_w_499);
AND_array_1509 AND_array_1509_i500(a,b[500],c_w_500);
AND_array_1509 AND_array_1509_i501(a,b[501],c_w_501);
AND_array_1509 AND_array_1509_i502(a,b[502],c_w_502);
AND_array_1509 AND_array_1509_i503(a,b[503],c_w_503);
AND_array_1509 AND_array_1509_i504(a,b[504],c_w_504);
AND_array_1509 AND_array_1509_i505(a,b[505],c_w_505);
AND_array_1509 AND_array_1509_i506(a,b[506],c_w_506);
AND_array_1509 AND_array_1509_i507(a,b[507],c_w_507);
AND_array_1509 AND_array_1509_i508(a,b[508],c_w_508);
AND_array_1509 AND_array_1509_i509(a,b[509],c_w_509);
AND_array_1509 AND_array_1509_i510(a,b[510],c_w_510);
AND_array_1509 AND_array_1509_i511(a,b[511],c_w_511);
AND_array_1509 AND_array_1509_i512(a,b[512],c_w_512);
AND_array_1509 AND_array_1509_i513(a,b[513],c_w_513);
AND_array_1509 AND_array_1509_i514(a,b[514],c_w_514);
AND_array_1509 AND_array_1509_i515(a,b[515],c_w_515);
AND_array_1509 AND_array_1509_i516(a,b[516],c_w_516);
AND_array_1509 AND_array_1509_i517(a,b[517],c_w_517);
AND_array_1509 AND_array_1509_i518(a,b[518],c_w_518);
AND_array_1509 AND_array_1509_i519(a,b[519],c_w_519);
AND_array_1509 AND_array_1509_i520(a,b[520],c_w_520);
AND_array_1509 AND_array_1509_i521(a,b[521],c_w_521);
AND_array_1509 AND_array_1509_i522(a,b[522],c_w_522);
AND_array_1509 AND_array_1509_i523(a,b[523],c_w_523);
AND_array_1509 AND_array_1509_i524(a,b[524],c_w_524);
AND_array_1509 AND_array_1509_i525(a,b[525],c_w_525);
AND_array_1509 AND_array_1509_i526(a,b[526],c_w_526);
AND_array_1509 AND_array_1509_i527(a,b[527],c_w_527);
AND_array_1509 AND_array_1509_i528(a,b[528],c_w_528);
AND_array_1509 AND_array_1509_i529(a,b[529],c_w_529);
AND_array_1509 AND_array_1509_i530(a,b[530],c_w_530);
AND_array_1509 AND_array_1509_i531(a,b[531],c_w_531);
AND_array_1509 AND_array_1509_i532(a,b[532],c_w_532);
AND_array_1509 AND_array_1509_i533(a,b[533],c_w_533);
AND_array_1509 AND_array_1509_i534(a,b[534],c_w_534);
AND_array_1509 AND_array_1509_i535(a,b[535],c_w_535);
AND_array_1509 AND_array_1509_i536(a,b[536],c_w_536);
AND_array_1509 AND_array_1509_i537(a,b[537],c_w_537);
AND_array_1509 AND_array_1509_i538(a,b[538],c_w_538);
AND_array_1509 AND_array_1509_i539(a,b[539],c_w_539);
AND_array_1509 AND_array_1509_i540(a,b[540],c_w_540);
AND_array_1509 AND_array_1509_i541(a,b[541],c_w_541);
AND_array_1509 AND_array_1509_i542(a,b[542],c_w_542);
AND_array_1509 AND_array_1509_i543(a,b[543],c_w_543);
AND_array_1509 AND_array_1509_i544(a,b[544],c_w_544);
AND_array_1509 AND_array_1509_i545(a,b[545],c_w_545);
AND_array_1509 AND_array_1509_i546(a,b[546],c_w_546);
AND_array_1509 AND_array_1509_i547(a,b[547],c_w_547);
AND_array_1509 AND_array_1509_i548(a,b[548],c_w_548);
AND_array_1509 AND_array_1509_i549(a,b[549],c_w_549);
AND_array_1509 AND_array_1509_i550(a,b[550],c_w_550);
AND_array_1509 AND_array_1509_i551(a,b[551],c_w_551);
AND_array_1509 AND_array_1509_i552(a,b[552],c_w_552);
AND_array_1509 AND_array_1509_i553(a,b[553],c_w_553);
AND_array_1509 AND_array_1509_i554(a,b[554],c_w_554);
AND_array_1509 AND_array_1509_i555(a,b[555],c_w_555);
AND_array_1509 AND_array_1509_i556(a,b[556],c_w_556);
AND_array_1509 AND_array_1509_i557(a,b[557],c_w_557);
AND_array_1509 AND_array_1509_i558(a,b[558],c_w_558);
AND_array_1509 AND_array_1509_i559(a,b[559],c_w_559);
AND_array_1509 AND_array_1509_i560(a,b[560],c_w_560);
AND_array_1509 AND_array_1509_i561(a,b[561],c_w_561);
AND_array_1509 AND_array_1509_i562(a,b[562],c_w_562);
AND_array_1509 AND_array_1509_i563(a,b[563],c_w_563);
AND_array_1509 AND_array_1509_i564(a,b[564],c_w_564);
AND_array_1509 AND_array_1509_i565(a,b[565],c_w_565);
AND_array_1509 AND_array_1509_i566(a,b[566],c_w_566);
AND_array_1509 AND_array_1509_i567(a,b[567],c_w_567);
AND_array_1509 AND_array_1509_i568(a,b[568],c_w_568);
AND_array_1509 AND_array_1509_i569(a,b[569],c_w_569);
AND_array_1509 AND_array_1509_i570(a,b[570],c_w_570);
AND_array_1509 AND_array_1509_i571(a,b[571],c_w_571);
AND_array_1509 AND_array_1509_i572(a,b[572],c_w_572);
AND_array_1509 AND_array_1509_i573(a,b[573],c_w_573);
AND_array_1509 AND_array_1509_i574(a,b[574],c_w_574);
AND_array_1509 AND_array_1509_i575(a,b[575],c_w_575);
AND_array_1509 AND_array_1509_i576(a,b[576],c_w_576);
AND_array_1509 AND_array_1509_i577(a,b[577],c_w_577);
AND_array_1509 AND_array_1509_i578(a,b[578],c_w_578);
AND_array_1509 AND_array_1509_i579(a,b[579],c_w_579);
AND_array_1509 AND_array_1509_i580(a,b[580],c_w_580);
AND_array_1509 AND_array_1509_i581(a,b[581],c_w_581);
AND_array_1509 AND_array_1509_i582(a,b[582],c_w_582);
AND_array_1509 AND_array_1509_i583(a,b[583],c_w_583);
AND_array_1509 AND_array_1509_i584(a,b[584],c_w_584);
AND_array_1509 AND_array_1509_i585(a,b[585],c_w_585);
AND_array_1509 AND_array_1509_i586(a,b[586],c_w_586);
AND_array_1509 AND_array_1509_i587(a,b[587],c_w_587);
AND_array_1509 AND_array_1509_i588(a,b[588],c_w_588);
AND_array_1509 AND_array_1509_i589(a,b[589],c_w_589);
AND_array_1509 AND_array_1509_i590(a,b[590],c_w_590);
AND_array_1509 AND_array_1509_i591(a,b[591],c_w_591);
AND_array_1509 AND_array_1509_i592(a,b[592],c_w_592);
AND_array_1509 AND_array_1509_i593(a,b[593],c_w_593);
AND_array_1509 AND_array_1509_i594(a,b[594],c_w_594);
AND_array_1509 AND_array_1509_i595(a,b[595],c_w_595);
AND_array_1509 AND_array_1509_i596(a,b[596],c_w_596);
AND_array_1509 AND_array_1509_i597(a,b[597],c_w_597);
AND_array_1509 AND_array_1509_i598(a,b[598],c_w_598);
AND_array_1509 AND_array_1509_i599(a,b[599],c_w_599);
AND_array_1509 AND_array_1509_i600(a,b[600],c_w_600);
AND_array_1509 AND_array_1509_i601(a,b[601],c_w_601);
AND_array_1509 AND_array_1509_i602(a,b[602],c_w_602);
AND_array_1509 AND_array_1509_i603(a,b[603],c_w_603);
AND_array_1509 AND_array_1509_i604(a,b[604],c_w_604);
AND_array_1509 AND_array_1509_i605(a,b[605],c_w_605);
AND_array_1509 AND_array_1509_i606(a,b[606],c_w_606);
AND_array_1509 AND_array_1509_i607(a,b[607],c_w_607);
AND_array_1509 AND_array_1509_i608(a,b[608],c_w_608);
AND_array_1509 AND_array_1509_i609(a,b[609],c_w_609);
AND_array_1509 AND_array_1509_i610(a,b[610],c_w_610);
AND_array_1509 AND_array_1509_i611(a,b[611],c_w_611);
AND_array_1509 AND_array_1509_i612(a,b[612],c_w_612);
AND_array_1509 AND_array_1509_i613(a,b[613],c_w_613);
AND_array_1509 AND_array_1509_i614(a,b[614],c_w_614);
AND_array_1509 AND_array_1509_i615(a,b[615],c_w_615);
AND_array_1509 AND_array_1509_i616(a,b[616],c_w_616);
AND_array_1509 AND_array_1509_i617(a,b[617],c_w_617);
AND_array_1509 AND_array_1509_i618(a,b[618],c_w_618);
AND_array_1509 AND_array_1509_i619(a,b[619],c_w_619);
AND_array_1509 AND_array_1509_i620(a,b[620],c_w_620);
AND_array_1509 AND_array_1509_i621(a,b[621],c_w_621);
AND_array_1509 AND_array_1509_i622(a,b[622],c_w_622);
AND_array_1509 AND_array_1509_i623(a,b[623],c_w_623);
AND_array_1509 AND_array_1509_i624(a,b[624],c_w_624);
AND_array_1509 AND_array_1509_i625(a,b[625],c_w_625);
AND_array_1509 AND_array_1509_i626(a,b[626],c_w_626);
AND_array_1509 AND_array_1509_i627(a,b[627],c_w_627);
AND_array_1509 AND_array_1509_i628(a,b[628],c_w_628);
AND_array_1509 AND_array_1509_i629(a,b[629],c_w_629);
AND_array_1509 AND_array_1509_i630(a,b[630],c_w_630);
AND_array_1509 AND_array_1509_i631(a,b[631],c_w_631);
AND_array_1509 AND_array_1509_i632(a,b[632],c_w_632);
AND_array_1509 AND_array_1509_i633(a,b[633],c_w_633);
AND_array_1509 AND_array_1509_i634(a,b[634],c_w_634);
AND_array_1509 AND_array_1509_i635(a,b[635],c_w_635);
AND_array_1509 AND_array_1509_i636(a,b[636],c_w_636);
AND_array_1509 AND_array_1509_i637(a,b[637],c_w_637);
AND_array_1509 AND_array_1509_i638(a,b[638],c_w_638);
AND_array_1509 AND_array_1509_i639(a,b[639],c_w_639);
AND_array_1509 AND_array_1509_i640(a,b[640],c_w_640);
AND_array_1509 AND_array_1509_i641(a,b[641],c_w_641);
AND_array_1509 AND_array_1509_i642(a,b[642],c_w_642);
AND_array_1509 AND_array_1509_i643(a,b[643],c_w_643);
AND_array_1509 AND_array_1509_i644(a,b[644],c_w_644);
AND_array_1509 AND_array_1509_i645(a,b[645],c_w_645);
AND_array_1509 AND_array_1509_i646(a,b[646],c_w_646);
AND_array_1509 AND_array_1509_i647(a,b[647],c_w_647);
AND_array_1509 AND_array_1509_i648(a,b[648],c_w_648);
AND_array_1509 AND_array_1509_i649(a,b[649],c_w_649);
AND_array_1509 AND_array_1509_i650(a,b[650],c_w_650);
AND_array_1509 AND_array_1509_i651(a,b[651],c_w_651);
AND_array_1509 AND_array_1509_i652(a,b[652],c_w_652);
AND_array_1509 AND_array_1509_i653(a,b[653],c_w_653);
AND_array_1509 AND_array_1509_i654(a,b[654],c_w_654);
AND_array_1509 AND_array_1509_i655(a,b[655],c_w_655);
AND_array_1509 AND_array_1509_i656(a,b[656],c_w_656);
AND_array_1509 AND_array_1509_i657(a,b[657],c_w_657);
AND_array_1509 AND_array_1509_i658(a,b[658],c_w_658);
AND_array_1509 AND_array_1509_i659(a,b[659],c_w_659);
AND_array_1509 AND_array_1509_i660(a,b[660],c_w_660);
AND_array_1509 AND_array_1509_i661(a,b[661],c_w_661);
AND_array_1509 AND_array_1509_i662(a,b[662],c_w_662);
AND_array_1509 AND_array_1509_i663(a,b[663],c_w_663);
AND_array_1509 AND_array_1509_i664(a,b[664],c_w_664);
AND_array_1509 AND_array_1509_i665(a,b[665],c_w_665);
AND_array_1509 AND_array_1509_i666(a,b[666],c_w_666);
AND_array_1509 AND_array_1509_i667(a,b[667],c_w_667);
AND_array_1509 AND_array_1509_i668(a,b[668],c_w_668);
AND_array_1509 AND_array_1509_i669(a,b[669],c_w_669);
AND_array_1509 AND_array_1509_i670(a,b[670],c_w_670);
AND_array_1509 AND_array_1509_i671(a,b[671],c_w_671);
AND_array_1509 AND_array_1509_i672(a,b[672],c_w_672);
AND_array_1509 AND_array_1509_i673(a,b[673],c_w_673);
AND_array_1509 AND_array_1509_i674(a,b[674],c_w_674);
AND_array_1509 AND_array_1509_i675(a,b[675],c_w_675);
AND_array_1509 AND_array_1509_i676(a,b[676],c_w_676);
AND_array_1509 AND_array_1509_i677(a,b[677],c_w_677);
AND_array_1509 AND_array_1509_i678(a,b[678],c_w_678);
AND_array_1509 AND_array_1509_i679(a,b[679],c_w_679);
AND_array_1509 AND_array_1509_i680(a,b[680],c_w_680);
AND_array_1509 AND_array_1509_i681(a,b[681],c_w_681);
AND_array_1509 AND_array_1509_i682(a,b[682],c_w_682);
AND_array_1509 AND_array_1509_i683(a,b[683],c_w_683);
AND_array_1509 AND_array_1509_i684(a,b[684],c_w_684);
AND_array_1509 AND_array_1509_i685(a,b[685],c_w_685);
AND_array_1509 AND_array_1509_i686(a,b[686],c_w_686);
AND_array_1509 AND_array_1509_i687(a,b[687],c_w_687);
AND_array_1509 AND_array_1509_i688(a,b[688],c_w_688);
AND_array_1509 AND_array_1509_i689(a,b[689],c_w_689);
AND_array_1509 AND_array_1509_i690(a,b[690],c_w_690);
AND_array_1509 AND_array_1509_i691(a,b[691],c_w_691);
AND_array_1509 AND_array_1509_i692(a,b[692],c_w_692);
AND_array_1509 AND_array_1509_i693(a,b[693],c_w_693);
AND_array_1509 AND_array_1509_i694(a,b[694],c_w_694);
AND_array_1509 AND_array_1509_i695(a,b[695],c_w_695);
AND_array_1509 AND_array_1509_i696(a,b[696],c_w_696);
AND_array_1509 AND_array_1509_i697(a,b[697],c_w_697);
AND_array_1509 AND_array_1509_i698(a,b[698],c_w_698);
AND_array_1509 AND_array_1509_i699(a,b[699],c_w_699);
AND_array_1509 AND_array_1509_i700(a,b[700],c_w_700);
AND_array_1509 AND_array_1509_i701(a,b[701],c_w_701);
AND_array_1509 AND_array_1509_i702(a,b[702],c_w_702);
AND_array_1509 AND_array_1509_i703(a,b[703],c_w_703);
AND_array_1509 AND_array_1509_i704(a,b[704],c_w_704);
AND_array_1509 AND_array_1509_i705(a,b[705],c_w_705);
AND_array_1509 AND_array_1509_i706(a,b[706],c_w_706);
AND_array_1509 AND_array_1509_i707(a,b[707],c_w_707);
AND_array_1509 AND_array_1509_i708(a,b[708],c_w_708);
AND_array_1509 AND_array_1509_i709(a,b[709],c_w_709);
AND_array_1509 AND_array_1509_i710(a,b[710],c_w_710);
AND_array_1509 AND_array_1509_i711(a,b[711],c_w_711);
AND_array_1509 AND_array_1509_i712(a,b[712],c_w_712);
AND_array_1509 AND_array_1509_i713(a,b[713],c_w_713);
AND_array_1509 AND_array_1509_i714(a,b[714],c_w_714);
AND_array_1509 AND_array_1509_i715(a,b[715],c_w_715);
AND_array_1509 AND_array_1509_i716(a,b[716],c_w_716);
AND_array_1509 AND_array_1509_i717(a,b[717],c_w_717);
AND_array_1509 AND_array_1509_i718(a,b[718],c_w_718);
AND_array_1509 AND_array_1509_i719(a,b[719],c_w_719);
AND_array_1509 AND_array_1509_i720(a,b[720],c_w_720);
AND_array_1509 AND_array_1509_i721(a,b[721],c_w_721);
AND_array_1509 AND_array_1509_i722(a,b[722],c_w_722);
AND_array_1509 AND_array_1509_i723(a,b[723],c_w_723);
AND_array_1509 AND_array_1509_i724(a,b[724],c_w_724);
AND_array_1509 AND_array_1509_i725(a,b[725],c_w_725);
AND_array_1509 AND_array_1509_i726(a,b[726],c_w_726);
AND_array_1509 AND_array_1509_i727(a,b[727],c_w_727);
AND_array_1509 AND_array_1509_i728(a,b[728],c_w_728);
AND_array_1509 AND_array_1509_i729(a,b[729],c_w_729);
AND_array_1509 AND_array_1509_i730(a,b[730],c_w_730);
AND_array_1509 AND_array_1509_i731(a,b[731],c_w_731);
AND_array_1509 AND_array_1509_i732(a,b[732],c_w_732);
AND_array_1509 AND_array_1509_i733(a,b[733],c_w_733);
AND_array_1509 AND_array_1509_i734(a,b[734],c_w_734);
AND_array_1509 AND_array_1509_i735(a,b[735],c_w_735);
AND_array_1509 AND_array_1509_i736(a,b[736],c_w_736);
AND_array_1509 AND_array_1509_i737(a,b[737],c_w_737);
AND_array_1509 AND_array_1509_i738(a,b[738],c_w_738);
AND_array_1509 AND_array_1509_i739(a,b[739],c_w_739);
AND_array_1509 AND_array_1509_i740(a,b[740],c_w_740);
AND_array_1509 AND_array_1509_i741(a,b[741],c_w_741);
AND_array_1509 AND_array_1509_i742(a,b[742],c_w_742);
AND_array_1509 AND_array_1509_i743(a,b[743],c_w_743);
AND_array_1509 AND_array_1509_i744(a,b[744],c_w_744);
AND_array_1509 AND_array_1509_i745(a,b[745],c_w_745);
AND_array_1509 AND_array_1509_i746(a,b[746],c_w_746);
AND_array_1509 AND_array_1509_i747(a,b[747],c_w_747);
AND_array_1509 AND_array_1509_i748(a,b[748],c_w_748);
AND_array_1509 AND_array_1509_i749(a,b[749],c_w_749);
AND_array_1509 AND_array_1509_i750(a,b[750],c_w_750);
AND_array_1509 AND_array_1509_i751(a,b[751],c_w_751);
AND_array_1509 AND_array_1509_i752(a,b[752],c_w_752);
AND_array_1509 AND_array_1509_i753(a,b[753],c_w_753);
AND_array_1509 AND_array_1509_i754(a,b[754],c_w_754);
AND_array_1509 AND_array_1509_i755(a,b[755],c_w_755);
AND_array_1509 AND_array_1509_i756(a,b[756],c_w_756);
AND_array_1509 AND_array_1509_i757(a,b[757],c_w_757);
AND_array_1509 AND_array_1509_i758(a,b[758],c_w_758);
AND_array_1509 AND_array_1509_i759(a,b[759],c_w_759);
AND_array_1509 AND_array_1509_i760(a,b[760],c_w_760);
AND_array_1509 AND_array_1509_i761(a,b[761],c_w_761);
AND_array_1509 AND_array_1509_i762(a,b[762],c_w_762);
AND_array_1509 AND_array_1509_i763(a,b[763],c_w_763);
AND_array_1509 AND_array_1509_i764(a,b[764],c_w_764);
AND_array_1509 AND_array_1509_i765(a,b[765],c_w_765);
AND_array_1509 AND_array_1509_i766(a,b[766],c_w_766);
AND_array_1509 AND_array_1509_i767(a,b[767],c_w_767);
AND_array_1509 AND_array_1509_i768(a,b[768],c_w_768);
AND_array_1509 AND_array_1509_i769(a,b[769],c_w_769);
AND_array_1509 AND_array_1509_i770(a,b[770],c_w_770);
AND_array_1509 AND_array_1509_i771(a,b[771],c_w_771);
AND_array_1509 AND_array_1509_i772(a,b[772],c_w_772);
AND_array_1509 AND_array_1509_i773(a,b[773],c_w_773);
AND_array_1509 AND_array_1509_i774(a,b[774],c_w_774);
AND_array_1509 AND_array_1509_i775(a,b[775],c_w_775);
AND_array_1509 AND_array_1509_i776(a,b[776],c_w_776);
AND_array_1509 AND_array_1509_i777(a,b[777],c_w_777);
AND_array_1509 AND_array_1509_i778(a,b[778],c_w_778);
AND_array_1509 AND_array_1509_i779(a,b[779],c_w_779);
AND_array_1509 AND_array_1509_i780(a,b[780],c_w_780);
AND_array_1509 AND_array_1509_i781(a,b[781],c_w_781);
AND_array_1509 AND_array_1509_i782(a,b[782],c_w_782);
AND_array_1509 AND_array_1509_i783(a,b[783],c_w_783);
AND_array_1509 AND_array_1509_i784(a,b[784],c_w_784);
AND_array_1509 AND_array_1509_i785(a,b[785],c_w_785);
AND_array_1509 AND_array_1509_i786(a,b[786],c_w_786);
AND_array_1509 AND_array_1509_i787(a,b[787],c_w_787);
AND_array_1509 AND_array_1509_i788(a,b[788],c_w_788);
AND_array_1509 AND_array_1509_i789(a,b[789],c_w_789);
AND_array_1509 AND_array_1509_i790(a,b[790],c_w_790);
AND_array_1509 AND_array_1509_i791(a,b[791],c_w_791);
AND_array_1509 AND_array_1509_i792(a,b[792],c_w_792);
AND_array_1509 AND_array_1509_i793(a,b[793],c_w_793);
AND_array_1509 AND_array_1509_i794(a,b[794],c_w_794);
AND_array_1509 AND_array_1509_i795(a,b[795],c_w_795);
AND_array_1509 AND_array_1509_i796(a,b[796],c_w_796);
AND_array_1509 AND_array_1509_i797(a,b[797],c_w_797);
AND_array_1509 AND_array_1509_i798(a,b[798],c_w_798);
AND_array_1509 AND_array_1509_i799(a,b[799],c_w_799);
AND_array_1509 AND_array_1509_i800(a,b[800],c_w_800);
AND_array_1509 AND_array_1509_i801(a,b[801],c_w_801);
AND_array_1509 AND_array_1509_i802(a,b[802],c_w_802);
AND_array_1509 AND_array_1509_i803(a,b[803],c_w_803);
AND_array_1509 AND_array_1509_i804(a,b[804],c_w_804);
AND_array_1509 AND_array_1509_i805(a,b[805],c_w_805);
AND_array_1509 AND_array_1509_i806(a,b[806],c_w_806);
AND_array_1509 AND_array_1509_i807(a,b[807],c_w_807);
AND_array_1509 AND_array_1509_i808(a,b[808],c_w_808);
AND_array_1509 AND_array_1509_i809(a,b[809],c_w_809);
AND_array_1509 AND_array_1509_i810(a,b[810],c_w_810);
AND_array_1509 AND_array_1509_i811(a,b[811],c_w_811);
AND_array_1509 AND_array_1509_i812(a,b[812],c_w_812);
AND_array_1509 AND_array_1509_i813(a,b[813],c_w_813);
AND_array_1509 AND_array_1509_i814(a,b[814],c_w_814);
AND_array_1509 AND_array_1509_i815(a,b[815],c_w_815);
AND_array_1509 AND_array_1509_i816(a,b[816],c_w_816);
AND_array_1509 AND_array_1509_i817(a,b[817],c_w_817);
AND_array_1509 AND_array_1509_i818(a,b[818],c_w_818);
AND_array_1509 AND_array_1509_i819(a,b[819],c_w_819);
AND_array_1509 AND_array_1509_i820(a,b[820],c_w_820);
AND_array_1509 AND_array_1509_i821(a,b[821],c_w_821);
AND_array_1509 AND_array_1509_i822(a,b[822],c_w_822);
AND_array_1509 AND_array_1509_i823(a,b[823],c_w_823);
AND_array_1509 AND_array_1509_i824(a,b[824],c_w_824);
AND_array_1509 AND_array_1509_i825(a,b[825],c_w_825);
AND_array_1509 AND_array_1509_i826(a,b[826],c_w_826);
AND_array_1509 AND_array_1509_i827(a,b[827],c_w_827);
AND_array_1509 AND_array_1509_i828(a,b[828],c_w_828);
AND_array_1509 AND_array_1509_i829(a,b[829],c_w_829);
AND_array_1509 AND_array_1509_i830(a,b[830],c_w_830);
AND_array_1509 AND_array_1509_i831(a,b[831],c_w_831);
AND_array_1509 AND_array_1509_i832(a,b[832],c_w_832);
AND_array_1509 AND_array_1509_i833(a,b[833],c_w_833);
AND_array_1509 AND_array_1509_i834(a,b[834],c_w_834);
AND_array_1509 AND_array_1509_i835(a,b[835],c_w_835);
AND_array_1509 AND_array_1509_i836(a,b[836],c_w_836);
AND_array_1509 AND_array_1509_i837(a,b[837],c_w_837);
AND_array_1509 AND_array_1509_i838(a,b[838],c_w_838);
AND_array_1509 AND_array_1509_i839(a,b[839],c_w_839);
AND_array_1509 AND_array_1509_i840(a,b[840],c_w_840);
AND_array_1509 AND_array_1509_i841(a,b[841],c_w_841);
AND_array_1509 AND_array_1509_i842(a,b[842],c_w_842);
AND_array_1509 AND_array_1509_i843(a,b[843],c_w_843);
AND_array_1509 AND_array_1509_i844(a,b[844],c_w_844);
AND_array_1509 AND_array_1509_i845(a,b[845],c_w_845);
AND_array_1509 AND_array_1509_i846(a,b[846],c_w_846);
AND_array_1509 AND_array_1509_i847(a,b[847],c_w_847);
AND_array_1509 AND_array_1509_i848(a,b[848],c_w_848);
AND_array_1509 AND_array_1509_i849(a,b[849],c_w_849);
AND_array_1509 AND_array_1509_i850(a,b[850],c_w_850);
AND_array_1509 AND_array_1509_i851(a,b[851],c_w_851);
AND_array_1509 AND_array_1509_i852(a,b[852],c_w_852);
AND_array_1509 AND_array_1509_i853(a,b[853],c_w_853);
AND_array_1509 AND_array_1509_i854(a,b[854],c_w_854);
AND_array_1509 AND_array_1509_i855(a,b[855],c_w_855);
AND_array_1509 AND_array_1509_i856(a,b[856],c_w_856);
AND_array_1509 AND_array_1509_i857(a,b[857],c_w_857);
AND_array_1509 AND_array_1509_i858(a,b[858],c_w_858);
AND_array_1509 AND_array_1509_i859(a,b[859],c_w_859);
AND_array_1509 AND_array_1509_i860(a,b[860],c_w_860);
AND_array_1509 AND_array_1509_i861(a,b[861],c_w_861);
AND_array_1509 AND_array_1509_i862(a,b[862],c_w_862);
AND_array_1509 AND_array_1509_i863(a,b[863],c_w_863);
AND_array_1509 AND_array_1509_i864(a,b[864],c_w_864);
AND_array_1509 AND_array_1509_i865(a,b[865],c_w_865);
AND_array_1509 AND_array_1509_i866(a,b[866],c_w_866);
AND_array_1509 AND_array_1509_i867(a,b[867],c_w_867);
AND_array_1509 AND_array_1509_i868(a,b[868],c_w_868);
AND_array_1509 AND_array_1509_i869(a,b[869],c_w_869);
AND_array_1509 AND_array_1509_i870(a,b[870],c_w_870);
AND_array_1509 AND_array_1509_i871(a,b[871],c_w_871);
AND_array_1509 AND_array_1509_i872(a,b[872],c_w_872);
AND_array_1509 AND_array_1509_i873(a,b[873],c_w_873);
AND_array_1509 AND_array_1509_i874(a,b[874],c_w_874);
AND_array_1509 AND_array_1509_i875(a,b[875],c_w_875);
AND_array_1509 AND_array_1509_i876(a,b[876],c_w_876);
AND_array_1509 AND_array_1509_i877(a,b[877],c_w_877);
AND_array_1509 AND_array_1509_i878(a,b[878],c_w_878);
AND_array_1509 AND_array_1509_i879(a,b[879],c_w_879);
AND_array_1509 AND_array_1509_i880(a,b[880],c_w_880);
AND_array_1509 AND_array_1509_i881(a,b[881],c_w_881);
AND_array_1509 AND_array_1509_i882(a,b[882],c_w_882);
AND_array_1509 AND_array_1509_i883(a,b[883],c_w_883);
AND_array_1509 AND_array_1509_i884(a,b[884],c_w_884);
AND_array_1509 AND_array_1509_i885(a,b[885],c_w_885);
AND_array_1509 AND_array_1509_i886(a,b[886],c_w_886);
AND_array_1509 AND_array_1509_i887(a,b[887],c_w_887);
AND_array_1509 AND_array_1509_i888(a,b[888],c_w_888);
AND_array_1509 AND_array_1509_i889(a,b[889],c_w_889);
AND_array_1509 AND_array_1509_i890(a,b[890],c_w_890);
AND_array_1509 AND_array_1509_i891(a,b[891],c_w_891);
AND_array_1509 AND_array_1509_i892(a,b[892],c_w_892);
AND_array_1509 AND_array_1509_i893(a,b[893],c_w_893);
AND_array_1509 AND_array_1509_i894(a,b[894],c_w_894);
AND_array_1509 AND_array_1509_i895(a,b[895],c_w_895);
AND_array_1509 AND_array_1509_i896(a,b[896],c_w_896);
AND_array_1509 AND_array_1509_i897(a,b[897],c_w_897);
AND_array_1509 AND_array_1509_i898(a,b[898],c_w_898);
AND_array_1509 AND_array_1509_i899(a,b[899],c_w_899);
AND_array_1509 AND_array_1509_i900(a,b[900],c_w_900);
AND_array_1509 AND_array_1509_i901(a,b[901],c_w_901);
AND_array_1509 AND_array_1509_i902(a,b[902],c_w_902);
AND_array_1509 AND_array_1509_i903(a,b[903],c_w_903);
AND_array_1509 AND_array_1509_i904(a,b[904],c_w_904);
AND_array_1509 AND_array_1509_i905(a,b[905],c_w_905);
AND_array_1509 AND_array_1509_i906(a,b[906],c_w_906);
AND_array_1509 AND_array_1509_i907(a,b[907],c_w_907);
AND_array_1509 AND_array_1509_i908(a,b[908],c_w_908);
AND_array_1509 AND_array_1509_i909(a,b[909],c_w_909);
AND_array_1509 AND_array_1509_i910(a,b[910],c_w_910);
AND_array_1509 AND_array_1509_i911(a,b[911],c_w_911);
AND_array_1509 AND_array_1509_i912(a,b[912],c_w_912);
AND_array_1509 AND_array_1509_i913(a,b[913],c_w_913);
AND_array_1509 AND_array_1509_i914(a,b[914],c_w_914);
AND_array_1509 AND_array_1509_i915(a,b[915],c_w_915);
AND_array_1509 AND_array_1509_i916(a,b[916],c_w_916);
AND_array_1509 AND_array_1509_i917(a,b[917],c_w_917);
AND_array_1509 AND_array_1509_i918(a,b[918],c_w_918);
AND_array_1509 AND_array_1509_i919(a,b[919],c_w_919);
AND_array_1509 AND_array_1509_i920(a,b[920],c_w_920);
AND_array_1509 AND_array_1509_i921(a,b[921],c_w_921);
AND_array_1509 AND_array_1509_i922(a,b[922],c_w_922);
AND_array_1509 AND_array_1509_i923(a,b[923],c_w_923);
AND_array_1509 AND_array_1509_i924(a,b[924],c_w_924);
AND_array_1509 AND_array_1509_i925(a,b[925],c_w_925);
AND_array_1509 AND_array_1509_i926(a,b[926],c_w_926);
AND_array_1509 AND_array_1509_i927(a,b[927],c_w_927);
AND_array_1509 AND_array_1509_i928(a,b[928],c_w_928);
AND_array_1509 AND_array_1509_i929(a,b[929],c_w_929);
AND_array_1509 AND_array_1509_i930(a,b[930],c_w_930);
AND_array_1509 AND_array_1509_i931(a,b[931],c_w_931);
AND_array_1509 AND_array_1509_i932(a,b[932],c_w_932);
AND_array_1509 AND_array_1509_i933(a,b[933],c_w_933);
AND_array_1509 AND_array_1509_i934(a,b[934],c_w_934);
AND_array_1509 AND_array_1509_i935(a,b[935],c_w_935);
AND_array_1509 AND_array_1509_i936(a,b[936],c_w_936);
AND_array_1509 AND_array_1509_i937(a,b[937],c_w_937);
AND_array_1509 AND_array_1509_i938(a,b[938],c_w_938);
AND_array_1509 AND_array_1509_i939(a,b[939],c_w_939);
AND_array_1509 AND_array_1509_i940(a,b[940],c_w_940);
AND_array_1509 AND_array_1509_i941(a,b[941],c_w_941);
AND_array_1509 AND_array_1509_i942(a,b[942],c_w_942);
AND_array_1509 AND_array_1509_i943(a,b[943],c_w_943);
AND_array_1509 AND_array_1509_i944(a,b[944],c_w_944);
AND_array_1509 AND_array_1509_i945(a,b[945],c_w_945);
AND_array_1509 AND_array_1509_i946(a,b[946],c_w_946);
AND_array_1509 AND_array_1509_i947(a,b[947],c_w_947);
AND_array_1509 AND_array_1509_i948(a,b[948],c_w_948);
AND_array_1509 AND_array_1509_i949(a,b[949],c_w_949);
AND_array_1509 AND_array_1509_i950(a,b[950],c_w_950);
AND_array_1509 AND_array_1509_i951(a,b[951],c_w_951);
AND_array_1509 AND_array_1509_i952(a,b[952],c_w_952);
AND_array_1509 AND_array_1509_i953(a,b[953],c_w_953);
AND_array_1509 AND_array_1509_i954(a,b[954],c_w_954);
AND_array_1509 AND_array_1509_i955(a,b[955],c_w_955);
AND_array_1509 AND_array_1509_i956(a,b[956],c_w_956);
AND_array_1509 AND_array_1509_i957(a,b[957],c_w_957);
AND_array_1509 AND_array_1509_i958(a,b[958],c_w_958);
AND_array_1509 AND_array_1509_i959(a,b[959],c_w_959);
AND_array_1509 AND_array_1509_i960(a,b[960],c_w_960);
AND_array_1509 AND_array_1509_i961(a,b[961],c_w_961);
AND_array_1509 AND_array_1509_i962(a,b[962],c_w_962);
AND_array_1509 AND_array_1509_i963(a,b[963],c_w_963);
AND_array_1509 AND_array_1509_i964(a,b[964],c_w_964);
AND_array_1509 AND_array_1509_i965(a,b[965],c_w_965);
AND_array_1509 AND_array_1509_i966(a,b[966],c_w_966);
AND_array_1509 AND_array_1509_i967(a,b[967],c_w_967);
AND_array_1509 AND_array_1509_i968(a,b[968],c_w_968);
AND_array_1509 AND_array_1509_i969(a,b[969],c_w_969);
AND_array_1509 AND_array_1509_i970(a,b[970],c_w_970);
AND_array_1509 AND_array_1509_i971(a,b[971],c_w_971);
AND_array_1509 AND_array_1509_i972(a,b[972],c_w_972);
AND_array_1509 AND_array_1509_i973(a,b[973],c_w_973);
AND_array_1509 AND_array_1509_i974(a,b[974],c_w_974);
AND_array_1509 AND_array_1509_i975(a,b[975],c_w_975);
AND_array_1509 AND_array_1509_i976(a,b[976],c_w_976);
AND_array_1509 AND_array_1509_i977(a,b[977],c_w_977);
AND_array_1509 AND_array_1509_i978(a,b[978],c_w_978);
AND_array_1509 AND_array_1509_i979(a,b[979],c_w_979);
AND_array_1509 AND_array_1509_i980(a,b[980],c_w_980);
AND_array_1509 AND_array_1509_i981(a,b[981],c_w_981);
AND_array_1509 AND_array_1509_i982(a,b[982],c_w_982);
AND_array_1509 AND_array_1509_i983(a,b[983],c_w_983);
AND_array_1509 AND_array_1509_i984(a,b[984],c_w_984);
AND_array_1509 AND_array_1509_i985(a,b[985],c_w_985);
AND_array_1509 AND_array_1509_i986(a,b[986],c_w_986);
AND_array_1509 AND_array_1509_i987(a,b[987],c_w_987);
AND_array_1509 AND_array_1509_i988(a,b[988],c_w_988);
AND_array_1509 AND_array_1509_i989(a,b[989],c_w_989);
AND_array_1509 AND_array_1509_i990(a,b[990],c_w_990);
AND_array_1509 AND_array_1509_i991(a,b[991],c_w_991);
AND_array_1509 AND_array_1509_i992(a,b[992],c_w_992);
AND_array_1509 AND_array_1509_i993(a,b[993],c_w_993);
AND_array_1509 AND_array_1509_i994(a,b[994],c_w_994);
AND_array_1509 AND_array_1509_i995(a,b[995],c_w_995);
AND_array_1509 AND_array_1509_i996(a,b[996],c_w_996);
AND_array_1509 AND_array_1509_i997(a,b[997],c_w_997);
AND_array_1509 AND_array_1509_i998(a,b[998],c_w_998);
AND_array_1509 AND_array_1509_i999(a,b[999],c_w_999);
AND_array_1509 AND_array_1509_i1000(a,b[1000],c_w_1000);
AND_array_1509 AND_array_1509_i1001(a,b[1001],c_w_1001);
AND_array_1509 AND_array_1509_i1002(a,b[1002],c_w_1002);
AND_array_1509 AND_array_1509_i1003(a,b[1003],c_w_1003);
AND_array_1509 AND_array_1509_i1004(a,b[1004],c_w_1004);
AND_array_1509 AND_array_1509_i1005(a,b[1005],c_w_1005);
AND_array_1509 AND_array_1509_i1006(a,b[1006],c_w_1006);
AND_array_1509 AND_array_1509_i1007(a,b[1007],c_w_1007);
AND_array_1509 AND_array_1509_i1008(a,b[1008],c_w_1008);
AND_array_1509 AND_array_1509_i1009(a,b[1009],c_w_1009);
AND_array_1509 AND_array_1509_i1010(a,b[1010],c_w_1010);
AND_array_1509 AND_array_1509_i1011(a,b[1011],c_w_1011);
AND_array_1509 AND_array_1509_i1012(a,b[1012],c_w_1012);
AND_array_1509 AND_array_1509_i1013(a,b[1013],c_w_1013);
AND_array_1509 AND_array_1509_i1014(a,b[1014],c_w_1014);
AND_array_1509 AND_array_1509_i1015(a,b[1015],c_w_1015);
AND_array_1509 AND_array_1509_i1016(a,b[1016],c_w_1016);
AND_array_1509 AND_array_1509_i1017(a,b[1017],c_w_1017);
AND_array_1509 AND_array_1509_i1018(a,b[1018],c_w_1018);
AND_array_1509 AND_array_1509_i1019(a,b[1019],c_w_1019);
AND_array_1509 AND_array_1509_i1020(a,b[1020],c_w_1020);
AND_array_1509 AND_array_1509_i1021(a,b[1021],c_w_1021);
AND_array_1509 AND_array_1509_i1022(a,b[1022],c_w_1022);
AND_array_1509 AND_array_1509_i1023(a,b[1023],c_w_1023);
AND_array_1509 AND_array_1509_i1024(a,b[1024],c_w_1024);
AND_array_1509 AND_array_1509_i1025(a,b[1025],c_w_1025);
AND_array_1509 AND_array_1509_i1026(a,b[1026],c_w_1026);
AND_array_1509 AND_array_1509_i1027(a,b[1027],c_w_1027);
AND_array_1509 AND_array_1509_i1028(a,b[1028],c_w_1028);
AND_array_1509 AND_array_1509_i1029(a,b[1029],c_w_1029);
AND_array_1509 AND_array_1509_i1030(a,b[1030],c_w_1030);
AND_array_1509 AND_array_1509_i1031(a,b[1031],c_w_1031);
AND_array_1509 AND_array_1509_i1032(a,b[1032],c_w_1032);
AND_array_1509 AND_array_1509_i1033(a,b[1033],c_w_1033);
AND_array_1509 AND_array_1509_i1034(a,b[1034],c_w_1034);
AND_array_1509 AND_array_1509_i1035(a,b[1035],c_w_1035);
AND_array_1509 AND_array_1509_i1036(a,b[1036],c_w_1036);
AND_array_1509 AND_array_1509_i1037(a,b[1037],c_w_1037);
AND_array_1509 AND_array_1509_i1038(a,b[1038],c_w_1038);
AND_array_1509 AND_array_1509_i1039(a,b[1039],c_w_1039);
AND_array_1509 AND_array_1509_i1040(a,b[1040],c_w_1040);
AND_array_1509 AND_array_1509_i1041(a,b[1041],c_w_1041);
AND_array_1509 AND_array_1509_i1042(a,b[1042],c_w_1042);
AND_array_1509 AND_array_1509_i1043(a,b[1043],c_w_1043);
AND_array_1509 AND_array_1509_i1044(a,b[1044],c_w_1044);
AND_array_1509 AND_array_1509_i1045(a,b[1045],c_w_1045);
AND_array_1509 AND_array_1509_i1046(a,b[1046],c_w_1046);
AND_array_1509 AND_array_1509_i1047(a,b[1047],c_w_1047);
AND_array_1509 AND_array_1509_i1048(a,b[1048],c_w_1048);
AND_array_1509 AND_array_1509_i1049(a,b[1049],c_w_1049);
AND_array_1509 AND_array_1509_i1050(a,b[1050],c_w_1050);
AND_array_1509 AND_array_1509_i1051(a,b[1051],c_w_1051);
AND_array_1509 AND_array_1509_i1052(a,b[1052],c_w_1052);
AND_array_1509 AND_array_1509_i1053(a,b[1053],c_w_1053);
AND_array_1509 AND_array_1509_i1054(a,b[1054],c_w_1054);
AND_array_1509 AND_array_1509_i1055(a,b[1055],c_w_1055);
AND_array_1509 AND_array_1509_i1056(a,b[1056],c_w_1056);
AND_array_1509 AND_array_1509_i1057(a,b[1057],c_w_1057);
AND_array_1509 AND_array_1509_i1058(a,b[1058],c_w_1058);
AND_array_1509 AND_array_1509_i1059(a,b[1059],c_w_1059);
AND_array_1509 AND_array_1509_i1060(a,b[1060],c_w_1060);
AND_array_1509 AND_array_1509_i1061(a,b[1061],c_w_1061);
AND_array_1509 AND_array_1509_i1062(a,b[1062],c_w_1062);
AND_array_1509 AND_array_1509_i1063(a,b[1063],c_w_1063);
AND_array_1509 AND_array_1509_i1064(a,b[1064],c_w_1064);
AND_array_1509 AND_array_1509_i1065(a,b[1065],c_w_1065);
AND_array_1509 AND_array_1509_i1066(a,b[1066],c_w_1066);
AND_array_1509 AND_array_1509_i1067(a,b[1067],c_w_1067);
AND_array_1509 AND_array_1509_i1068(a,b[1068],c_w_1068);
AND_array_1509 AND_array_1509_i1069(a,b[1069],c_w_1069);
AND_array_1509 AND_array_1509_i1070(a,b[1070],c_w_1070);
AND_array_1509 AND_array_1509_i1071(a,b[1071],c_w_1071);
AND_array_1509 AND_array_1509_i1072(a,b[1072],c_w_1072);
AND_array_1509 AND_array_1509_i1073(a,b[1073],c_w_1073);
AND_array_1509 AND_array_1509_i1074(a,b[1074],c_w_1074);
AND_array_1509 AND_array_1509_i1075(a,b[1075],c_w_1075);
AND_array_1509 AND_array_1509_i1076(a,b[1076],c_w_1076);
AND_array_1509 AND_array_1509_i1077(a,b[1077],c_w_1077);
AND_array_1509 AND_array_1509_i1078(a,b[1078],c_w_1078);
AND_array_1509 AND_array_1509_i1079(a,b[1079],c_w_1079);
AND_array_1509 AND_array_1509_i1080(a,b[1080],c_w_1080);
AND_array_1509 AND_array_1509_i1081(a,b[1081],c_w_1081);
AND_array_1509 AND_array_1509_i1082(a,b[1082],c_w_1082);
AND_array_1509 AND_array_1509_i1083(a,b[1083],c_w_1083);
AND_array_1509 AND_array_1509_i1084(a,b[1084],c_w_1084);
AND_array_1509 AND_array_1509_i1085(a,b[1085],c_w_1085);
AND_array_1509 AND_array_1509_i1086(a,b[1086],c_w_1086);
AND_array_1509 AND_array_1509_i1087(a,b[1087],c_w_1087);
AND_array_1509 AND_array_1509_i1088(a,b[1088],c_w_1088);
AND_array_1509 AND_array_1509_i1089(a,b[1089],c_w_1089);
AND_array_1509 AND_array_1509_i1090(a,b[1090],c_w_1090);
AND_array_1509 AND_array_1509_i1091(a,b[1091],c_w_1091);
AND_array_1509 AND_array_1509_i1092(a,b[1092],c_w_1092);
AND_array_1509 AND_array_1509_i1093(a,b[1093],c_w_1093);
AND_array_1509 AND_array_1509_i1094(a,b[1094],c_w_1094);
AND_array_1509 AND_array_1509_i1095(a,b[1095],c_w_1095);
AND_array_1509 AND_array_1509_i1096(a,b[1096],c_w_1096);
AND_array_1509 AND_array_1509_i1097(a,b[1097],c_w_1097);
AND_array_1509 AND_array_1509_i1098(a,b[1098],c_w_1098);
AND_array_1509 AND_array_1509_i1099(a,b[1099],c_w_1099);
AND_array_1509 AND_array_1509_i1100(a,b[1100],c_w_1100);
AND_array_1509 AND_array_1509_i1101(a,b[1101],c_w_1101);
AND_array_1509 AND_array_1509_i1102(a,b[1102],c_w_1102);
AND_array_1509 AND_array_1509_i1103(a,b[1103],c_w_1103);
AND_array_1509 AND_array_1509_i1104(a,b[1104],c_w_1104);
AND_array_1509 AND_array_1509_i1105(a,b[1105],c_w_1105);
AND_array_1509 AND_array_1509_i1106(a,b[1106],c_w_1106);
AND_array_1509 AND_array_1509_i1107(a,b[1107],c_w_1107);
AND_array_1509 AND_array_1509_i1108(a,b[1108],c_w_1108);
AND_array_1509 AND_array_1509_i1109(a,b[1109],c_w_1109);
AND_array_1509 AND_array_1509_i1110(a,b[1110],c_w_1110);
AND_array_1509 AND_array_1509_i1111(a,b[1111],c_w_1111);
AND_array_1509 AND_array_1509_i1112(a,b[1112],c_w_1112);
AND_array_1509 AND_array_1509_i1113(a,b[1113],c_w_1113);
AND_array_1509 AND_array_1509_i1114(a,b[1114],c_w_1114);
AND_array_1509 AND_array_1509_i1115(a,b[1115],c_w_1115);
AND_array_1509 AND_array_1509_i1116(a,b[1116],c_w_1116);
AND_array_1509 AND_array_1509_i1117(a,b[1117],c_w_1117);
AND_array_1509 AND_array_1509_i1118(a,b[1118],c_w_1118);
AND_array_1509 AND_array_1509_i1119(a,b[1119],c_w_1119);
AND_array_1509 AND_array_1509_i1120(a,b[1120],c_w_1120);
AND_array_1509 AND_array_1509_i1121(a,b[1121],c_w_1121);
AND_array_1509 AND_array_1509_i1122(a,b[1122],c_w_1122);
AND_array_1509 AND_array_1509_i1123(a,b[1123],c_w_1123);
AND_array_1509 AND_array_1509_i1124(a,b[1124],c_w_1124);
AND_array_1509 AND_array_1509_i1125(a,b[1125],c_w_1125);
AND_array_1509 AND_array_1509_i1126(a,b[1126],c_w_1126);
AND_array_1509 AND_array_1509_i1127(a,b[1127],c_w_1127);
AND_array_1509 AND_array_1509_i1128(a,b[1128],c_w_1128);
AND_array_1509 AND_array_1509_i1129(a,b[1129],c_w_1129);
AND_array_1509 AND_array_1509_i1130(a,b[1130],c_w_1130);
AND_array_1509 AND_array_1509_i1131(a,b[1131],c_w_1131);
AND_array_1509 AND_array_1509_i1132(a,b[1132],c_w_1132);
AND_array_1509 AND_array_1509_i1133(a,b[1133],c_w_1133);
AND_array_1509 AND_array_1509_i1134(a,b[1134],c_w_1134);
AND_array_1509 AND_array_1509_i1135(a,b[1135],c_w_1135);
AND_array_1509 AND_array_1509_i1136(a,b[1136],c_w_1136);
AND_array_1509 AND_array_1509_i1137(a,b[1137],c_w_1137);
AND_array_1509 AND_array_1509_i1138(a,b[1138],c_w_1138);
AND_array_1509 AND_array_1509_i1139(a,b[1139],c_w_1139);
AND_array_1509 AND_array_1509_i1140(a,b[1140],c_w_1140);
AND_array_1509 AND_array_1509_i1141(a,b[1141],c_w_1141);
AND_array_1509 AND_array_1509_i1142(a,b[1142],c_w_1142);
AND_array_1509 AND_array_1509_i1143(a,b[1143],c_w_1143);
AND_array_1509 AND_array_1509_i1144(a,b[1144],c_w_1144);
AND_array_1509 AND_array_1509_i1145(a,b[1145],c_w_1145);
AND_array_1509 AND_array_1509_i1146(a,b[1146],c_w_1146);
AND_array_1509 AND_array_1509_i1147(a,b[1147],c_w_1147);
AND_array_1509 AND_array_1509_i1148(a,b[1148],c_w_1148);
AND_array_1509 AND_array_1509_i1149(a,b[1149],c_w_1149);
AND_array_1509 AND_array_1509_i1150(a,b[1150],c_w_1150);
AND_array_1509 AND_array_1509_i1151(a,b[1151],c_w_1151);
AND_array_1509 AND_array_1509_i1152(a,b[1152],c_w_1152);
AND_array_1509 AND_array_1509_i1153(a,b[1153],c_w_1153);
AND_array_1509 AND_array_1509_i1154(a,b[1154],c_w_1154);
AND_array_1509 AND_array_1509_i1155(a,b[1155],c_w_1155);
AND_array_1509 AND_array_1509_i1156(a,b[1156],c_w_1156);
AND_array_1509 AND_array_1509_i1157(a,b[1157],c_w_1157);
AND_array_1509 AND_array_1509_i1158(a,b[1158],c_w_1158);
AND_array_1509 AND_array_1509_i1159(a,b[1159],c_w_1159);
AND_array_1509 AND_array_1509_i1160(a,b[1160],c_w_1160);
AND_array_1509 AND_array_1509_i1161(a,b[1161],c_w_1161);
AND_array_1509 AND_array_1509_i1162(a,b[1162],c_w_1162);
AND_array_1509 AND_array_1509_i1163(a,b[1163],c_w_1163);
AND_array_1509 AND_array_1509_i1164(a,b[1164],c_w_1164);
AND_array_1509 AND_array_1509_i1165(a,b[1165],c_w_1165);
AND_array_1509 AND_array_1509_i1166(a,b[1166],c_w_1166);
AND_array_1509 AND_array_1509_i1167(a,b[1167],c_w_1167);
AND_array_1509 AND_array_1509_i1168(a,b[1168],c_w_1168);
AND_array_1509 AND_array_1509_i1169(a,b[1169],c_w_1169);
AND_array_1509 AND_array_1509_i1170(a,b[1170],c_w_1170);
AND_array_1509 AND_array_1509_i1171(a,b[1171],c_w_1171);
AND_array_1509 AND_array_1509_i1172(a,b[1172],c_w_1172);
AND_array_1509 AND_array_1509_i1173(a,b[1173],c_w_1173);
AND_array_1509 AND_array_1509_i1174(a,b[1174],c_w_1174);
AND_array_1509 AND_array_1509_i1175(a,b[1175],c_w_1175);
AND_array_1509 AND_array_1509_i1176(a,b[1176],c_w_1176);
AND_array_1509 AND_array_1509_i1177(a,b[1177],c_w_1177);
AND_array_1509 AND_array_1509_i1178(a,b[1178],c_w_1178);
AND_array_1509 AND_array_1509_i1179(a,b[1179],c_w_1179);
AND_array_1509 AND_array_1509_i1180(a,b[1180],c_w_1180);
AND_array_1509 AND_array_1509_i1181(a,b[1181],c_w_1181);
AND_array_1509 AND_array_1509_i1182(a,b[1182],c_w_1182);
AND_array_1509 AND_array_1509_i1183(a,b[1183],c_w_1183);
AND_array_1509 AND_array_1509_i1184(a,b[1184],c_w_1184);
AND_array_1509 AND_array_1509_i1185(a,b[1185],c_w_1185);
AND_array_1509 AND_array_1509_i1186(a,b[1186],c_w_1186);
AND_array_1509 AND_array_1509_i1187(a,b[1187],c_w_1187);
AND_array_1509 AND_array_1509_i1188(a,b[1188],c_w_1188);
AND_array_1509 AND_array_1509_i1189(a,b[1189],c_w_1189);
AND_array_1509 AND_array_1509_i1190(a,b[1190],c_w_1190);
AND_array_1509 AND_array_1509_i1191(a,b[1191],c_w_1191);
AND_array_1509 AND_array_1509_i1192(a,b[1192],c_w_1192);
AND_array_1509 AND_array_1509_i1193(a,b[1193],c_w_1193);
AND_array_1509 AND_array_1509_i1194(a,b[1194],c_w_1194);
AND_array_1509 AND_array_1509_i1195(a,b[1195],c_w_1195);
AND_array_1509 AND_array_1509_i1196(a,b[1196],c_w_1196);
AND_array_1509 AND_array_1509_i1197(a,b[1197],c_w_1197);
AND_array_1509 AND_array_1509_i1198(a,b[1198],c_w_1198);
AND_array_1509 AND_array_1509_i1199(a,b[1199],c_w_1199);
AND_array_1509 AND_array_1509_i1200(a,b[1200],c_w_1200);
AND_array_1509 AND_array_1509_i1201(a,b[1201],c_w_1201);
AND_array_1509 AND_array_1509_i1202(a,b[1202],c_w_1202);
AND_array_1509 AND_array_1509_i1203(a,b[1203],c_w_1203);
AND_array_1509 AND_array_1509_i1204(a,b[1204],c_w_1204);
AND_array_1509 AND_array_1509_i1205(a,b[1205],c_w_1205);
AND_array_1509 AND_array_1509_i1206(a,b[1206],c_w_1206);
AND_array_1509 AND_array_1509_i1207(a,b[1207],c_w_1207);
AND_array_1509 AND_array_1509_i1208(a,b[1208],c_w_1208);
AND_array_1509 AND_array_1509_i1209(a,b[1209],c_w_1209);
AND_array_1509 AND_array_1509_i1210(a,b[1210],c_w_1210);
AND_array_1509 AND_array_1509_i1211(a,b[1211],c_w_1211);
AND_array_1509 AND_array_1509_i1212(a,b[1212],c_w_1212);
AND_array_1509 AND_array_1509_i1213(a,b[1213],c_w_1213);
AND_array_1509 AND_array_1509_i1214(a,b[1214],c_w_1214);
AND_array_1509 AND_array_1509_i1215(a,b[1215],c_w_1215);
AND_array_1509 AND_array_1509_i1216(a,b[1216],c_w_1216);
AND_array_1509 AND_array_1509_i1217(a,b[1217],c_w_1217);
AND_array_1509 AND_array_1509_i1218(a,b[1218],c_w_1218);
AND_array_1509 AND_array_1509_i1219(a,b[1219],c_w_1219);
AND_array_1509 AND_array_1509_i1220(a,b[1220],c_w_1220);
AND_array_1509 AND_array_1509_i1221(a,b[1221],c_w_1221);
AND_array_1509 AND_array_1509_i1222(a,b[1222],c_w_1222);
AND_array_1509 AND_array_1509_i1223(a,b[1223],c_w_1223);
AND_array_1509 AND_array_1509_i1224(a,b[1224],c_w_1224);
AND_array_1509 AND_array_1509_i1225(a,b[1225],c_w_1225);
AND_array_1509 AND_array_1509_i1226(a,b[1226],c_w_1226);
AND_array_1509 AND_array_1509_i1227(a,b[1227],c_w_1227);
AND_array_1509 AND_array_1509_i1228(a,b[1228],c_w_1228);
AND_array_1509 AND_array_1509_i1229(a,b[1229],c_w_1229);
AND_array_1509 AND_array_1509_i1230(a,b[1230],c_w_1230);
AND_array_1509 AND_array_1509_i1231(a,b[1231],c_w_1231);
AND_array_1509 AND_array_1509_i1232(a,b[1232],c_w_1232);
AND_array_1509 AND_array_1509_i1233(a,b[1233],c_w_1233);
AND_array_1509 AND_array_1509_i1234(a,b[1234],c_w_1234);
AND_array_1509 AND_array_1509_i1235(a,b[1235],c_w_1235);
AND_array_1509 AND_array_1509_i1236(a,b[1236],c_w_1236);
AND_array_1509 AND_array_1509_i1237(a,b[1237],c_w_1237);
AND_array_1509 AND_array_1509_i1238(a,b[1238],c_w_1238);
AND_array_1509 AND_array_1509_i1239(a,b[1239],c_w_1239);
AND_array_1509 AND_array_1509_i1240(a,b[1240],c_w_1240);
AND_array_1509 AND_array_1509_i1241(a,b[1241],c_w_1241);
AND_array_1509 AND_array_1509_i1242(a,b[1242],c_w_1242);
AND_array_1509 AND_array_1509_i1243(a,b[1243],c_w_1243);
AND_array_1509 AND_array_1509_i1244(a,b[1244],c_w_1244);
AND_array_1509 AND_array_1509_i1245(a,b[1245],c_w_1245);
AND_array_1509 AND_array_1509_i1246(a,b[1246],c_w_1246);
AND_array_1509 AND_array_1509_i1247(a,b[1247],c_w_1247);
AND_array_1509 AND_array_1509_i1248(a,b[1248],c_w_1248);
AND_array_1509 AND_array_1509_i1249(a,b[1249],c_w_1249);
AND_array_1509 AND_array_1509_i1250(a,b[1250],c_w_1250);
AND_array_1509 AND_array_1509_i1251(a,b[1251],c_w_1251);
AND_array_1509 AND_array_1509_i1252(a,b[1252],c_w_1252);
AND_array_1509 AND_array_1509_i1253(a,b[1253],c_w_1253);
AND_array_1509 AND_array_1509_i1254(a,b[1254],c_w_1254);
AND_array_1509 AND_array_1509_i1255(a,b[1255],c_w_1255);
AND_array_1509 AND_array_1509_i1256(a,b[1256],c_w_1256);
AND_array_1509 AND_array_1509_i1257(a,b[1257],c_w_1257);
AND_array_1509 AND_array_1509_i1258(a,b[1258],c_w_1258);
AND_array_1509 AND_array_1509_i1259(a,b[1259],c_w_1259);
AND_array_1509 AND_array_1509_i1260(a,b[1260],c_w_1260);
AND_array_1509 AND_array_1509_i1261(a,b[1261],c_w_1261);
AND_array_1509 AND_array_1509_i1262(a,b[1262],c_w_1262);
AND_array_1509 AND_array_1509_i1263(a,b[1263],c_w_1263);
AND_array_1509 AND_array_1509_i1264(a,b[1264],c_w_1264);
AND_array_1509 AND_array_1509_i1265(a,b[1265],c_w_1265);
AND_array_1509 AND_array_1509_i1266(a,b[1266],c_w_1266);
AND_array_1509 AND_array_1509_i1267(a,b[1267],c_w_1267);
AND_array_1509 AND_array_1509_i1268(a,b[1268],c_w_1268);
AND_array_1509 AND_array_1509_i1269(a,b[1269],c_w_1269);
AND_array_1509 AND_array_1509_i1270(a,b[1270],c_w_1270);
AND_array_1509 AND_array_1509_i1271(a,b[1271],c_w_1271);
AND_array_1509 AND_array_1509_i1272(a,b[1272],c_w_1272);
AND_array_1509 AND_array_1509_i1273(a,b[1273],c_w_1273);
AND_array_1509 AND_array_1509_i1274(a,b[1274],c_w_1274);
AND_array_1509 AND_array_1509_i1275(a,b[1275],c_w_1275);
AND_array_1509 AND_array_1509_i1276(a,b[1276],c_w_1276);
AND_array_1509 AND_array_1509_i1277(a,b[1277],c_w_1277);
AND_array_1509 AND_array_1509_i1278(a,b[1278],c_w_1278);
AND_array_1509 AND_array_1509_i1279(a,b[1279],c_w_1279);
AND_array_1509 AND_array_1509_i1280(a,b[1280],c_w_1280);
AND_array_1509 AND_array_1509_i1281(a,b[1281],c_w_1281);
AND_array_1509 AND_array_1509_i1282(a,b[1282],c_w_1282);
AND_array_1509 AND_array_1509_i1283(a,b[1283],c_w_1283);
AND_array_1509 AND_array_1509_i1284(a,b[1284],c_w_1284);
AND_array_1509 AND_array_1509_i1285(a,b[1285],c_w_1285);
AND_array_1509 AND_array_1509_i1286(a,b[1286],c_w_1286);
AND_array_1509 AND_array_1509_i1287(a,b[1287],c_w_1287);
AND_array_1509 AND_array_1509_i1288(a,b[1288],c_w_1288);
AND_array_1509 AND_array_1509_i1289(a,b[1289],c_w_1289);
AND_array_1509 AND_array_1509_i1290(a,b[1290],c_w_1290);
AND_array_1509 AND_array_1509_i1291(a,b[1291],c_w_1291);
AND_array_1509 AND_array_1509_i1292(a,b[1292],c_w_1292);
AND_array_1509 AND_array_1509_i1293(a,b[1293],c_w_1293);
AND_array_1509 AND_array_1509_i1294(a,b[1294],c_w_1294);
AND_array_1509 AND_array_1509_i1295(a,b[1295],c_w_1295);
AND_array_1509 AND_array_1509_i1296(a,b[1296],c_w_1296);
AND_array_1509 AND_array_1509_i1297(a,b[1297],c_w_1297);
AND_array_1509 AND_array_1509_i1298(a,b[1298],c_w_1298);
AND_array_1509 AND_array_1509_i1299(a,b[1299],c_w_1299);
AND_array_1509 AND_array_1509_i1300(a,b[1300],c_w_1300);
AND_array_1509 AND_array_1509_i1301(a,b[1301],c_w_1301);
AND_array_1509 AND_array_1509_i1302(a,b[1302],c_w_1302);
AND_array_1509 AND_array_1509_i1303(a,b[1303],c_w_1303);
AND_array_1509 AND_array_1509_i1304(a,b[1304],c_w_1304);
AND_array_1509 AND_array_1509_i1305(a,b[1305],c_w_1305);
AND_array_1509 AND_array_1509_i1306(a,b[1306],c_w_1306);
AND_array_1509 AND_array_1509_i1307(a,b[1307],c_w_1307);
AND_array_1509 AND_array_1509_i1308(a,b[1308],c_w_1308);
AND_array_1509 AND_array_1509_i1309(a,b[1309],c_w_1309);
AND_array_1509 AND_array_1509_i1310(a,b[1310],c_w_1310);
AND_array_1509 AND_array_1509_i1311(a,b[1311],c_w_1311);
AND_array_1509 AND_array_1509_i1312(a,b[1312],c_w_1312);
AND_array_1509 AND_array_1509_i1313(a,b[1313],c_w_1313);
AND_array_1509 AND_array_1509_i1314(a,b[1314],c_w_1314);
AND_array_1509 AND_array_1509_i1315(a,b[1315],c_w_1315);
AND_array_1509 AND_array_1509_i1316(a,b[1316],c_w_1316);
AND_array_1509 AND_array_1509_i1317(a,b[1317],c_w_1317);
AND_array_1509 AND_array_1509_i1318(a,b[1318],c_w_1318);
AND_array_1509 AND_array_1509_i1319(a,b[1319],c_w_1319);
AND_array_1509 AND_array_1509_i1320(a,b[1320],c_w_1320);
AND_array_1509 AND_array_1509_i1321(a,b[1321],c_w_1321);
AND_array_1509 AND_array_1509_i1322(a,b[1322],c_w_1322);
AND_array_1509 AND_array_1509_i1323(a,b[1323],c_w_1323);
AND_array_1509 AND_array_1509_i1324(a,b[1324],c_w_1324);
AND_array_1509 AND_array_1509_i1325(a,b[1325],c_w_1325);
AND_array_1509 AND_array_1509_i1326(a,b[1326],c_w_1326);
AND_array_1509 AND_array_1509_i1327(a,b[1327],c_w_1327);
AND_array_1509 AND_array_1509_i1328(a,b[1328],c_w_1328);
AND_array_1509 AND_array_1509_i1329(a,b[1329],c_w_1329);
AND_array_1509 AND_array_1509_i1330(a,b[1330],c_w_1330);
AND_array_1509 AND_array_1509_i1331(a,b[1331],c_w_1331);
AND_array_1509 AND_array_1509_i1332(a,b[1332],c_w_1332);
AND_array_1509 AND_array_1509_i1333(a,b[1333],c_w_1333);
AND_array_1509 AND_array_1509_i1334(a,b[1334],c_w_1334);
AND_array_1509 AND_array_1509_i1335(a,b[1335],c_w_1335);
AND_array_1509 AND_array_1509_i1336(a,b[1336],c_w_1336);
AND_array_1509 AND_array_1509_i1337(a,b[1337],c_w_1337);
AND_array_1509 AND_array_1509_i1338(a,b[1338],c_w_1338);
AND_array_1509 AND_array_1509_i1339(a,b[1339],c_w_1339);
AND_array_1509 AND_array_1509_i1340(a,b[1340],c_w_1340);
AND_array_1509 AND_array_1509_i1341(a,b[1341],c_w_1341);
AND_array_1509 AND_array_1509_i1342(a,b[1342],c_w_1342);
AND_array_1509 AND_array_1509_i1343(a,b[1343],c_w_1343);
AND_array_1509 AND_array_1509_i1344(a,b[1344],c_w_1344);
AND_array_1509 AND_array_1509_i1345(a,b[1345],c_w_1345);
AND_array_1509 AND_array_1509_i1346(a,b[1346],c_w_1346);
AND_array_1509 AND_array_1509_i1347(a,b[1347],c_w_1347);
AND_array_1509 AND_array_1509_i1348(a,b[1348],c_w_1348);
AND_array_1509 AND_array_1509_i1349(a,b[1349],c_w_1349);
AND_array_1509 AND_array_1509_i1350(a,b[1350],c_w_1350);
AND_array_1509 AND_array_1509_i1351(a,b[1351],c_w_1351);
AND_array_1509 AND_array_1509_i1352(a,b[1352],c_w_1352);
AND_array_1509 AND_array_1509_i1353(a,b[1353],c_w_1353);
AND_array_1509 AND_array_1509_i1354(a,b[1354],c_w_1354);
AND_array_1509 AND_array_1509_i1355(a,b[1355],c_w_1355);
AND_array_1509 AND_array_1509_i1356(a,b[1356],c_w_1356);
AND_array_1509 AND_array_1509_i1357(a,b[1357],c_w_1357);
AND_array_1509 AND_array_1509_i1358(a,b[1358],c_w_1358);
AND_array_1509 AND_array_1509_i1359(a,b[1359],c_w_1359);
AND_array_1509 AND_array_1509_i1360(a,b[1360],c_w_1360);
AND_array_1509 AND_array_1509_i1361(a,b[1361],c_w_1361);
AND_array_1509 AND_array_1509_i1362(a,b[1362],c_w_1362);
AND_array_1509 AND_array_1509_i1363(a,b[1363],c_w_1363);
AND_array_1509 AND_array_1509_i1364(a,b[1364],c_w_1364);
AND_array_1509 AND_array_1509_i1365(a,b[1365],c_w_1365);
AND_array_1509 AND_array_1509_i1366(a,b[1366],c_w_1366);
AND_array_1509 AND_array_1509_i1367(a,b[1367],c_w_1367);
AND_array_1509 AND_array_1509_i1368(a,b[1368],c_w_1368);
AND_array_1509 AND_array_1509_i1369(a,b[1369],c_w_1369);
AND_array_1509 AND_array_1509_i1370(a,b[1370],c_w_1370);
AND_array_1509 AND_array_1509_i1371(a,b[1371],c_w_1371);
AND_array_1509 AND_array_1509_i1372(a,b[1372],c_w_1372);
AND_array_1509 AND_array_1509_i1373(a,b[1373],c_w_1373);
AND_array_1509 AND_array_1509_i1374(a,b[1374],c_w_1374);
AND_array_1509 AND_array_1509_i1375(a,b[1375],c_w_1375);
AND_array_1509 AND_array_1509_i1376(a,b[1376],c_w_1376);
AND_array_1509 AND_array_1509_i1377(a,b[1377],c_w_1377);
AND_array_1509 AND_array_1509_i1378(a,b[1378],c_w_1378);
AND_array_1509 AND_array_1509_i1379(a,b[1379],c_w_1379);
AND_array_1509 AND_array_1509_i1380(a,b[1380],c_w_1380);
AND_array_1509 AND_array_1509_i1381(a,b[1381],c_w_1381);
AND_array_1509 AND_array_1509_i1382(a,b[1382],c_w_1382);
AND_array_1509 AND_array_1509_i1383(a,b[1383],c_w_1383);
AND_array_1509 AND_array_1509_i1384(a,b[1384],c_w_1384);
AND_array_1509 AND_array_1509_i1385(a,b[1385],c_w_1385);
AND_array_1509 AND_array_1509_i1386(a,b[1386],c_w_1386);
AND_array_1509 AND_array_1509_i1387(a,b[1387],c_w_1387);
AND_array_1509 AND_array_1509_i1388(a,b[1388],c_w_1388);
AND_array_1509 AND_array_1509_i1389(a,b[1389],c_w_1389);
AND_array_1509 AND_array_1509_i1390(a,b[1390],c_w_1390);
AND_array_1509 AND_array_1509_i1391(a,b[1391],c_w_1391);
AND_array_1509 AND_array_1509_i1392(a,b[1392],c_w_1392);
AND_array_1509 AND_array_1509_i1393(a,b[1393],c_w_1393);
AND_array_1509 AND_array_1509_i1394(a,b[1394],c_w_1394);
AND_array_1509 AND_array_1509_i1395(a,b[1395],c_w_1395);
AND_array_1509 AND_array_1509_i1396(a,b[1396],c_w_1396);
AND_array_1509 AND_array_1509_i1397(a,b[1397],c_w_1397);
AND_array_1509 AND_array_1509_i1398(a,b[1398],c_w_1398);
AND_array_1509 AND_array_1509_i1399(a,b[1399],c_w_1399);
AND_array_1509 AND_array_1509_i1400(a,b[1400],c_w_1400);
AND_array_1509 AND_array_1509_i1401(a,b[1401],c_w_1401);
AND_array_1509 AND_array_1509_i1402(a,b[1402],c_w_1402);
AND_array_1509 AND_array_1509_i1403(a,b[1403],c_w_1403);
AND_array_1509 AND_array_1509_i1404(a,b[1404],c_w_1404);
AND_array_1509 AND_array_1509_i1405(a,b[1405],c_w_1405);
AND_array_1509 AND_array_1509_i1406(a,b[1406],c_w_1406);
AND_array_1509 AND_array_1509_i1407(a,b[1407],c_w_1407);
AND_array_1509 AND_array_1509_i1408(a,b[1408],c_w_1408);
AND_array_1509 AND_array_1509_i1409(a,b[1409],c_w_1409);
AND_array_1509 AND_array_1509_i1410(a,b[1410],c_w_1410);
AND_array_1509 AND_array_1509_i1411(a,b[1411],c_w_1411);
AND_array_1509 AND_array_1509_i1412(a,b[1412],c_w_1412);
AND_array_1509 AND_array_1509_i1413(a,b[1413],c_w_1413);
AND_array_1509 AND_array_1509_i1414(a,b[1414],c_w_1414);
AND_array_1509 AND_array_1509_i1415(a,b[1415],c_w_1415);
AND_array_1509 AND_array_1509_i1416(a,b[1416],c_w_1416);
AND_array_1509 AND_array_1509_i1417(a,b[1417],c_w_1417);
AND_array_1509 AND_array_1509_i1418(a,b[1418],c_w_1418);
AND_array_1509 AND_array_1509_i1419(a,b[1419],c_w_1419);
AND_array_1509 AND_array_1509_i1420(a,b[1420],c_w_1420);
AND_array_1509 AND_array_1509_i1421(a,b[1421],c_w_1421);
AND_array_1509 AND_array_1509_i1422(a,b[1422],c_w_1422);
AND_array_1509 AND_array_1509_i1423(a,b[1423],c_w_1423);
AND_array_1509 AND_array_1509_i1424(a,b[1424],c_w_1424);
AND_array_1509 AND_array_1509_i1425(a,b[1425],c_w_1425);
AND_array_1509 AND_array_1509_i1426(a,b[1426],c_w_1426);
AND_array_1509 AND_array_1509_i1427(a,b[1427],c_w_1427);
AND_array_1509 AND_array_1509_i1428(a,b[1428],c_w_1428);
AND_array_1509 AND_array_1509_i1429(a,b[1429],c_w_1429);
AND_array_1509 AND_array_1509_i1430(a,b[1430],c_w_1430);
AND_array_1509 AND_array_1509_i1431(a,b[1431],c_w_1431);
AND_array_1509 AND_array_1509_i1432(a,b[1432],c_w_1432);
AND_array_1509 AND_array_1509_i1433(a,b[1433],c_w_1433);
AND_array_1509 AND_array_1509_i1434(a,b[1434],c_w_1434);
AND_array_1509 AND_array_1509_i1435(a,b[1435],c_w_1435);
AND_array_1509 AND_array_1509_i1436(a,b[1436],c_w_1436);
AND_array_1509 AND_array_1509_i1437(a,b[1437],c_w_1437);
AND_array_1509 AND_array_1509_i1438(a,b[1438],c_w_1438);
AND_array_1509 AND_array_1509_i1439(a,b[1439],c_w_1439);
AND_array_1509 AND_array_1509_i1440(a,b[1440],c_w_1440);
AND_array_1509 AND_array_1509_i1441(a,b[1441],c_w_1441);
AND_array_1509 AND_array_1509_i1442(a,b[1442],c_w_1442);
AND_array_1509 AND_array_1509_i1443(a,b[1443],c_w_1443);
AND_array_1509 AND_array_1509_i1444(a,b[1444],c_w_1444);
AND_array_1509 AND_array_1509_i1445(a,b[1445],c_w_1445);
AND_array_1509 AND_array_1509_i1446(a,b[1446],c_w_1446);
AND_array_1509 AND_array_1509_i1447(a,b[1447],c_w_1447);
AND_array_1509 AND_array_1509_i1448(a,b[1448],c_w_1448);
AND_array_1509 AND_array_1509_i1449(a,b[1449],c_w_1449);
AND_array_1509 AND_array_1509_i1450(a,b[1450],c_w_1450);
AND_array_1509 AND_array_1509_i1451(a,b[1451],c_w_1451);
AND_array_1509 AND_array_1509_i1452(a,b[1452],c_w_1452);
AND_array_1509 AND_array_1509_i1453(a,b[1453],c_w_1453);
AND_array_1509 AND_array_1509_i1454(a,b[1454],c_w_1454);
AND_array_1509 AND_array_1509_i1455(a,b[1455],c_w_1455);
AND_array_1509 AND_array_1509_i1456(a,b[1456],c_w_1456);
AND_array_1509 AND_array_1509_i1457(a,b[1457],c_w_1457);
AND_array_1509 AND_array_1509_i1458(a,b[1458],c_w_1458);
AND_array_1509 AND_array_1509_i1459(a,b[1459],c_w_1459);
AND_array_1509 AND_array_1509_i1460(a,b[1460],c_w_1460);
AND_array_1509 AND_array_1509_i1461(a,b[1461],c_w_1461);
AND_array_1509 AND_array_1509_i1462(a,b[1462],c_w_1462);
AND_array_1509 AND_array_1509_i1463(a,b[1463],c_w_1463);
AND_array_1509 AND_array_1509_i1464(a,b[1464],c_w_1464);
AND_array_1509 AND_array_1509_i1465(a,b[1465],c_w_1465);
AND_array_1509 AND_array_1509_i1466(a,b[1466],c_w_1466);
AND_array_1509 AND_array_1509_i1467(a,b[1467],c_w_1467);
AND_array_1509 AND_array_1509_i1468(a,b[1468],c_w_1468);
AND_array_1509 AND_array_1509_i1469(a,b[1469],c_w_1469);
AND_array_1509 AND_array_1509_i1470(a,b[1470],c_w_1470);
AND_array_1509 AND_array_1509_i1471(a,b[1471],c_w_1471);
AND_array_1509 AND_array_1509_i1472(a,b[1472],c_w_1472);
AND_array_1509 AND_array_1509_i1473(a,b[1473],c_w_1473);
AND_array_1509 AND_array_1509_i1474(a,b[1474],c_w_1474);
AND_array_1509 AND_array_1509_i1475(a,b[1475],c_w_1475);
AND_array_1509 AND_array_1509_i1476(a,b[1476],c_w_1476);
AND_array_1509 AND_array_1509_i1477(a,b[1477],c_w_1477);
AND_array_1509 AND_array_1509_i1478(a,b[1478],c_w_1478);
AND_array_1509 AND_array_1509_i1479(a,b[1479],c_w_1479);
AND_array_1509 AND_array_1509_i1480(a,b[1480],c_w_1480);
AND_array_1509 AND_array_1509_i1481(a,b[1481],c_w_1481);
AND_array_1509 AND_array_1509_i1482(a,b[1482],c_w_1482);
AND_array_1509 AND_array_1509_i1483(a,b[1483],c_w_1483);
AND_array_1509 AND_array_1509_i1484(a,b[1484],c_w_1484);
AND_array_1509 AND_array_1509_i1485(a,b[1485],c_w_1485);
AND_array_1509 AND_array_1509_i1486(a,b[1486],c_w_1486);
AND_array_1509 AND_array_1509_i1487(a,b[1487],c_w_1487);
AND_array_1509 AND_array_1509_i1488(a,b[1488],c_w_1488);
AND_array_1509 AND_array_1509_i1489(a,b[1489],c_w_1489);
AND_array_1509 AND_array_1509_i1490(a,b[1490],c_w_1490);
AND_array_1509 AND_array_1509_i1491(a,b[1491],c_w_1491);
AND_array_1509 AND_array_1509_i1492(a,b[1492],c_w_1492);
AND_array_1509 AND_array_1509_i1493(a,b[1493],c_w_1493);
AND_array_1509 AND_array_1509_i1494(a,b[1494],c_w_1494);
AND_array_1509 AND_array_1509_i1495(a,b[1495],c_w_1495);
AND_array_1509 AND_array_1509_i1496(a,b[1496],c_w_1496);
AND_array_1509 AND_array_1509_i1497(a,b[1497],c_w_1497);
AND_array_1509 AND_array_1509_i1498(a,b[1498],c_w_1498);
AND_array_1509 AND_array_1509_i1499(a,b[1499],c_w_1499);
AND_array_1509 AND_array_1509_i1500(a,b[1500],c_w_1500);
AND_array_1509 AND_array_1509_i1501(a,b[1501],c_w_1501);
AND_array_1509 AND_array_1509_i1502(a,b[1502],c_w_1502);
AND_array_1509 AND_array_1509_i1503(a,b[1503],c_w_1503);
AND_array_1509 AND_array_1509_i1504(a,b[1504],c_w_1504);
AND_array_1509 AND_array_1509_i1505(a,b[1505],c_w_1505);
AND_array_1509 AND_array_1509_i1506(a,b[1506],c_w_1506);
AND_array_1509 AND_array_1509_i1507(a,b[1507],c_w_1507);
AND_array_1509 AND_array_1509_i1508(a,b[1508],c_w_1508);
    
assign c[3017:0] = {1509'b0,c_w_0};
assign c[6035:3018] = {1508'b0,c_w_1,1'b0};
assign c[9053:6036] = {1507'b0,c_w_2,2'b0};
assign c[12071:9054] = {1506'b0,c_w_3,3'b0};
assign c[15089:12072] = {1505'b0,c_w_4,4'b0};
assign c[18107:15090] = {1504'b0,c_w_5,5'b0};
assign c[21125:18108] = {1503'b0,c_w_6,6'b0};
assign c[24143:21126] = {1502'b0,c_w_7,7'b0};
assign c[27161:24144] = {1501'b0,c_w_8,8'b0};
assign c[30179:27162] = {1500'b0,c_w_9,9'b0};
assign c[33197:30180] = {1499'b0,c_w_10,10'b0};
assign c[36215:33198] = {1498'b0,c_w_11,11'b0};
assign c[39233:36216] = {1497'b0,c_w_12,12'b0};
assign c[42251:39234] = {1496'b0,c_w_13,13'b0};
assign c[45269:42252] = {1495'b0,c_w_14,14'b0};
assign c[48287:45270] = {1494'b0,c_w_15,15'b0};
assign c[51305:48288] = {1493'b0,c_w_16,16'b0};
assign c[54323:51306] = {1492'b0,c_w_17,17'b0};
assign c[57341:54324] = {1491'b0,c_w_18,18'b0};
assign c[60359:57342] = {1490'b0,c_w_19,19'b0};
assign c[63377:60360] = {1489'b0,c_w_20,20'b0};
assign c[66395:63378] = {1488'b0,c_w_21,21'b0};
assign c[69413:66396] = {1487'b0,c_w_22,22'b0};
assign c[72431:69414] = {1486'b0,c_w_23,23'b0};
assign c[75449:72432] = {1485'b0,c_w_24,24'b0};
assign c[78467:75450] = {1484'b0,c_w_25,25'b0};
assign c[81485:78468] = {1483'b0,c_w_26,26'b0};
assign c[84503:81486] = {1482'b0,c_w_27,27'b0};
assign c[87521:84504] = {1481'b0,c_w_28,28'b0};
assign c[90539:87522] = {1480'b0,c_w_29,29'b0};
assign c[93557:90540] = {1479'b0,c_w_30,30'b0};
assign c[96575:93558] = {1478'b0,c_w_31,31'b0};
assign c[99593:96576] = {1477'b0,c_w_32,32'b0};
assign c[102611:99594] = {1476'b0,c_w_33,33'b0};
assign c[105629:102612] = {1475'b0,c_w_34,34'b0};
assign c[108647:105630] = {1474'b0,c_w_35,35'b0};
assign c[111665:108648] = {1473'b0,c_w_36,36'b0};
assign c[114683:111666] = {1472'b0,c_w_37,37'b0};
assign c[117701:114684] = {1471'b0,c_w_38,38'b0};
assign c[120719:117702] = {1470'b0,c_w_39,39'b0};
assign c[123737:120720] = {1469'b0,c_w_40,40'b0};
assign c[126755:123738] = {1468'b0,c_w_41,41'b0};
assign c[129773:126756] = {1467'b0,c_w_42,42'b0};
assign c[132791:129774] = {1466'b0,c_w_43,43'b0};
assign c[135809:132792] = {1465'b0,c_w_44,44'b0};
assign c[138827:135810] = {1464'b0,c_w_45,45'b0};
assign c[141845:138828] = {1463'b0,c_w_46,46'b0};
assign c[144863:141846] = {1462'b0,c_w_47,47'b0};
assign c[147881:144864] = {1461'b0,c_w_48,48'b0};
assign c[150899:147882] = {1460'b0,c_w_49,49'b0};
assign c[153917:150900] = {1459'b0,c_w_50,50'b0};
assign c[156935:153918] = {1458'b0,c_w_51,51'b0};
assign c[159953:156936] = {1457'b0,c_w_52,52'b0};
assign c[162971:159954] = {1456'b0,c_w_53,53'b0};
assign c[165989:162972] = {1455'b0,c_w_54,54'b0};
assign c[169007:165990] = {1454'b0,c_w_55,55'b0};
assign c[172025:169008] = {1453'b0,c_w_56,56'b0};
assign c[175043:172026] = {1452'b0,c_w_57,57'b0};
assign c[178061:175044] = {1451'b0,c_w_58,58'b0};
assign c[181079:178062] = {1450'b0,c_w_59,59'b0};
assign c[184097:181080] = {1449'b0,c_w_60,60'b0};
assign c[187115:184098] = {1448'b0,c_w_61,61'b0};
assign c[190133:187116] = {1447'b0,c_w_62,62'b0};
assign c[193151:190134] = {1446'b0,c_w_63,63'b0};
assign c[196169:193152] = {1445'b0,c_w_64,64'b0};
assign c[199187:196170] = {1444'b0,c_w_65,65'b0};
assign c[202205:199188] = {1443'b0,c_w_66,66'b0};
assign c[205223:202206] = {1442'b0,c_w_67,67'b0};
assign c[208241:205224] = {1441'b0,c_w_68,68'b0};
assign c[211259:208242] = {1440'b0,c_w_69,69'b0};
assign c[214277:211260] = {1439'b0,c_w_70,70'b0};
assign c[217295:214278] = {1438'b0,c_w_71,71'b0};
assign c[220313:217296] = {1437'b0,c_w_72,72'b0};
assign c[223331:220314] = {1436'b0,c_w_73,73'b0};
assign c[226349:223332] = {1435'b0,c_w_74,74'b0};
assign c[229367:226350] = {1434'b0,c_w_75,75'b0};
assign c[232385:229368] = {1433'b0,c_w_76,76'b0};
assign c[235403:232386] = {1432'b0,c_w_77,77'b0};
assign c[238421:235404] = {1431'b0,c_w_78,78'b0};
assign c[241439:238422] = {1430'b0,c_w_79,79'b0};
assign c[244457:241440] = {1429'b0,c_w_80,80'b0};
assign c[247475:244458] = {1428'b0,c_w_81,81'b0};
assign c[250493:247476] = {1427'b0,c_w_82,82'b0};
assign c[253511:250494] = {1426'b0,c_w_83,83'b0};
assign c[256529:253512] = {1425'b0,c_w_84,84'b0};
assign c[259547:256530] = {1424'b0,c_w_85,85'b0};
assign c[262565:259548] = {1423'b0,c_w_86,86'b0};
assign c[265583:262566] = {1422'b0,c_w_87,87'b0};
assign c[268601:265584] = {1421'b0,c_w_88,88'b0};
assign c[271619:268602] = {1420'b0,c_w_89,89'b0};
assign c[274637:271620] = {1419'b0,c_w_90,90'b0};
assign c[277655:274638] = {1418'b0,c_w_91,91'b0};
assign c[280673:277656] = {1417'b0,c_w_92,92'b0};
assign c[283691:280674] = {1416'b0,c_w_93,93'b0};
assign c[286709:283692] = {1415'b0,c_w_94,94'b0};
assign c[289727:286710] = {1414'b0,c_w_95,95'b0};
assign c[292745:289728] = {1413'b0,c_w_96,96'b0};
assign c[295763:292746] = {1412'b0,c_w_97,97'b0};
assign c[298781:295764] = {1411'b0,c_w_98,98'b0};
assign c[301799:298782] = {1410'b0,c_w_99,99'b0};
assign c[304817:301800] = {1409'b0,c_w_100,100'b0};
assign c[307835:304818] = {1408'b0,c_w_101,101'b0};
assign c[310853:307836] = {1407'b0,c_w_102,102'b0};
assign c[313871:310854] = {1406'b0,c_w_103,103'b0};
assign c[316889:313872] = {1405'b0,c_w_104,104'b0};
assign c[319907:316890] = {1404'b0,c_w_105,105'b0};
assign c[322925:319908] = {1403'b0,c_w_106,106'b0};
assign c[325943:322926] = {1402'b0,c_w_107,107'b0};
assign c[328961:325944] = {1401'b0,c_w_108,108'b0};
assign c[331979:328962] = {1400'b0,c_w_109,109'b0};
assign c[334997:331980] = {1399'b0,c_w_110,110'b0};
assign c[338015:334998] = {1398'b0,c_w_111,111'b0};
assign c[341033:338016] = {1397'b0,c_w_112,112'b0};
assign c[344051:341034] = {1396'b0,c_w_113,113'b0};
assign c[347069:344052] = {1395'b0,c_w_114,114'b0};
assign c[350087:347070] = {1394'b0,c_w_115,115'b0};
assign c[353105:350088] = {1393'b0,c_w_116,116'b0};
assign c[356123:353106] = {1392'b0,c_w_117,117'b0};
assign c[359141:356124] = {1391'b0,c_w_118,118'b0};
assign c[362159:359142] = {1390'b0,c_w_119,119'b0};
assign c[365177:362160] = {1389'b0,c_w_120,120'b0};
assign c[368195:365178] = {1388'b0,c_w_121,121'b0};
assign c[371213:368196] = {1387'b0,c_w_122,122'b0};
assign c[374231:371214] = {1386'b0,c_w_123,123'b0};
assign c[377249:374232] = {1385'b0,c_w_124,124'b0};
assign c[380267:377250] = {1384'b0,c_w_125,125'b0};
assign c[383285:380268] = {1383'b0,c_w_126,126'b0};
assign c[386303:383286] = {1382'b0,c_w_127,127'b0};
assign c[389321:386304] = {1381'b0,c_w_128,128'b0};
assign c[392339:389322] = {1380'b0,c_w_129,129'b0};
assign c[395357:392340] = {1379'b0,c_w_130,130'b0};
assign c[398375:395358] = {1378'b0,c_w_131,131'b0};
assign c[401393:398376] = {1377'b0,c_w_132,132'b0};
assign c[404411:401394] = {1376'b0,c_w_133,133'b0};
assign c[407429:404412] = {1375'b0,c_w_134,134'b0};
assign c[410447:407430] = {1374'b0,c_w_135,135'b0};
assign c[413465:410448] = {1373'b0,c_w_136,136'b0};
assign c[416483:413466] = {1372'b0,c_w_137,137'b0};
assign c[419501:416484] = {1371'b0,c_w_138,138'b0};
assign c[422519:419502] = {1370'b0,c_w_139,139'b0};
assign c[425537:422520] = {1369'b0,c_w_140,140'b0};
assign c[428555:425538] = {1368'b0,c_w_141,141'b0};
assign c[431573:428556] = {1367'b0,c_w_142,142'b0};
assign c[434591:431574] = {1366'b0,c_w_143,143'b0};
assign c[437609:434592] = {1365'b0,c_w_144,144'b0};
assign c[440627:437610] = {1364'b0,c_w_145,145'b0};
assign c[443645:440628] = {1363'b0,c_w_146,146'b0};
assign c[446663:443646] = {1362'b0,c_w_147,147'b0};
assign c[449681:446664] = {1361'b0,c_w_148,148'b0};
assign c[452699:449682] = {1360'b0,c_w_149,149'b0};
assign c[455717:452700] = {1359'b0,c_w_150,150'b0};
assign c[458735:455718] = {1358'b0,c_w_151,151'b0};
assign c[461753:458736] = {1357'b0,c_w_152,152'b0};
assign c[464771:461754] = {1356'b0,c_w_153,153'b0};
assign c[467789:464772] = {1355'b0,c_w_154,154'b0};
assign c[470807:467790] = {1354'b0,c_w_155,155'b0};
assign c[473825:470808] = {1353'b0,c_w_156,156'b0};
assign c[476843:473826] = {1352'b0,c_w_157,157'b0};
assign c[479861:476844] = {1351'b0,c_w_158,158'b0};
assign c[482879:479862] = {1350'b0,c_w_159,159'b0};
assign c[485897:482880] = {1349'b0,c_w_160,160'b0};
assign c[488915:485898] = {1348'b0,c_w_161,161'b0};
assign c[491933:488916] = {1347'b0,c_w_162,162'b0};
assign c[494951:491934] = {1346'b0,c_w_163,163'b0};
assign c[497969:494952] = {1345'b0,c_w_164,164'b0};
assign c[500987:497970] = {1344'b0,c_w_165,165'b0};
assign c[504005:500988] = {1343'b0,c_w_166,166'b0};
assign c[507023:504006] = {1342'b0,c_w_167,167'b0};
assign c[510041:507024] = {1341'b0,c_w_168,168'b0};
assign c[513059:510042] = {1340'b0,c_w_169,169'b0};
assign c[516077:513060] = {1339'b0,c_w_170,170'b0};
assign c[519095:516078] = {1338'b0,c_w_171,171'b0};
assign c[522113:519096] = {1337'b0,c_w_172,172'b0};
assign c[525131:522114] = {1336'b0,c_w_173,173'b0};
assign c[528149:525132] = {1335'b0,c_w_174,174'b0};
assign c[531167:528150] = {1334'b0,c_w_175,175'b0};
assign c[534185:531168] = {1333'b0,c_w_176,176'b0};
assign c[537203:534186] = {1332'b0,c_w_177,177'b0};
assign c[540221:537204] = {1331'b0,c_w_178,178'b0};
assign c[543239:540222] = {1330'b0,c_w_179,179'b0};
assign c[546257:543240] = {1329'b0,c_w_180,180'b0};
assign c[549275:546258] = {1328'b0,c_w_181,181'b0};
assign c[552293:549276] = {1327'b0,c_w_182,182'b0};
assign c[555311:552294] = {1326'b0,c_w_183,183'b0};
assign c[558329:555312] = {1325'b0,c_w_184,184'b0};
assign c[561347:558330] = {1324'b0,c_w_185,185'b0};
assign c[564365:561348] = {1323'b0,c_w_186,186'b0};
assign c[567383:564366] = {1322'b0,c_w_187,187'b0};
assign c[570401:567384] = {1321'b0,c_w_188,188'b0};
assign c[573419:570402] = {1320'b0,c_w_189,189'b0};
assign c[576437:573420] = {1319'b0,c_w_190,190'b0};
assign c[579455:576438] = {1318'b0,c_w_191,191'b0};
assign c[582473:579456] = {1317'b0,c_w_192,192'b0};
assign c[585491:582474] = {1316'b0,c_w_193,193'b0};
assign c[588509:585492] = {1315'b0,c_w_194,194'b0};
assign c[591527:588510] = {1314'b0,c_w_195,195'b0};
assign c[594545:591528] = {1313'b0,c_w_196,196'b0};
assign c[597563:594546] = {1312'b0,c_w_197,197'b0};
assign c[600581:597564] = {1311'b0,c_w_198,198'b0};
assign c[603599:600582] = {1310'b0,c_w_199,199'b0};
assign c[606617:603600] = {1309'b0,c_w_200,200'b0};
assign c[609635:606618] = {1308'b0,c_w_201,201'b0};
assign c[612653:609636] = {1307'b0,c_w_202,202'b0};
assign c[615671:612654] = {1306'b0,c_w_203,203'b0};
assign c[618689:615672] = {1305'b0,c_w_204,204'b0};
assign c[621707:618690] = {1304'b0,c_w_205,205'b0};
assign c[624725:621708] = {1303'b0,c_w_206,206'b0};
assign c[627743:624726] = {1302'b0,c_w_207,207'b0};
assign c[630761:627744] = {1301'b0,c_w_208,208'b0};
assign c[633779:630762] = {1300'b0,c_w_209,209'b0};
assign c[636797:633780] = {1299'b0,c_w_210,210'b0};
assign c[639815:636798] = {1298'b0,c_w_211,211'b0};
assign c[642833:639816] = {1297'b0,c_w_212,212'b0};
assign c[645851:642834] = {1296'b0,c_w_213,213'b0};
assign c[648869:645852] = {1295'b0,c_w_214,214'b0};
assign c[651887:648870] = {1294'b0,c_w_215,215'b0};
assign c[654905:651888] = {1293'b0,c_w_216,216'b0};
assign c[657923:654906] = {1292'b0,c_w_217,217'b0};
assign c[660941:657924] = {1291'b0,c_w_218,218'b0};
assign c[663959:660942] = {1290'b0,c_w_219,219'b0};
assign c[666977:663960] = {1289'b0,c_w_220,220'b0};
assign c[669995:666978] = {1288'b0,c_w_221,221'b0};
assign c[673013:669996] = {1287'b0,c_w_222,222'b0};
assign c[676031:673014] = {1286'b0,c_w_223,223'b0};
assign c[679049:676032] = {1285'b0,c_w_224,224'b0};
assign c[682067:679050] = {1284'b0,c_w_225,225'b0};
assign c[685085:682068] = {1283'b0,c_w_226,226'b0};
assign c[688103:685086] = {1282'b0,c_w_227,227'b0};
assign c[691121:688104] = {1281'b0,c_w_228,228'b0};
assign c[694139:691122] = {1280'b0,c_w_229,229'b0};
assign c[697157:694140] = {1279'b0,c_w_230,230'b0};
assign c[700175:697158] = {1278'b0,c_w_231,231'b0};
assign c[703193:700176] = {1277'b0,c_w_232,232'b0};
assign c[706211:703194] = {1276'b0,c_w_233,233'b0};
assign c[709229:706212] = {1275'b0,c_w_234,234'b0};
assign c[712247:709230] = {1274'b0,c_w_235,235'b0};
assign c[715265:712248] = {1273'b0,c_w_236,236'b0};
assign c[718283:715266] = {1272'b0,c_w_237,237'b0};
assign c[721301:718284] = {1271'b0,c_w_238,238'b0};
assign c[724319:721302] = {1270'b0,c_w_239,239'b0};
assign c[727337:724320] = {1269'b0,c_w_240,240'b0};
assign c[730355:727338] = {1268'b0,c_w_241,241'b0};
assign c[733373:730356] = {1267'b0,c_w_242,242'b0};
assign c[736391:733374] = {1266'b0,c_w_243,243'b0};
assign c[739409:736392] = {1265'b0,c_w_244,244'b0};
assign c[742427:739410] = {1264'b0,c_w_245,245'b0};
assign c[745445:742428] = {1263'b0,c_w_246,246'b0};
assign c[748463:745446] = {1262'b0,c_w_247,247'b0};
assign c[751481:748464] = {1261'b0,c_w_248,248'b0};
assign c[754499:751482] = {1260'b0,c_w_249,249'b0};
assign c[757517:754500] = {1259'b0,c_w_250,250'b0};
assign c[760535:757518] = {1258'b0,c_w_251,251'b0};
assign c[763553:760536] = {1257'b0,c_w_252,252'b0};
assign c[766571:763554] = {1256'b0,c_w_253,253'b0};
assign c[769589:766572] = {1255'b0,c_w_254,254'b0};
assign c[772607:769590] = {1254'b0,c_w_255,255'b0};
assign c[775625:772608] = {1253'b0,c_w_256,256'b0};
assign c[778643:775626] = {1252'b0,c_w_257,257'b0};
assign c[781661:778644] = {1251'b0,c_w_258,258'b0};
assign c[784679:781662] = {1250'b0,c_w_259,259'b0};
assign c[787697:784680] = {1249'b0,c_w_260,260'b0};
assign c[790715:787698] = {1248'b0,c_w_261,261'b0};
assign c[793733:790716] = {1247'b0,c_w_262,262'b0};
assign c[796751:793734] = {1246'b0,c_w_263,263'b0};
assign c[799769:796752] = {1245'b0,c_w_264,264'b0};
assign c[802787:799770] = {1244'b0,c_w_265,265'b0};
assign c[805805:802788] = {1243'b0,c_w_266,266'b0};
assign c[808823:805806] = {1242'b0,c_w_267,267'b0};
assign c[811841:808824] = {1241'b0,c_w_268,268'b0};
assign c[814859:811842] = {1240'b0,c_w_269,269'b0};
assign c[817877:814860] = {1239'b0,c_w_270,270'b0};
assign c[820895:817878] = {1238'b0,c_w_271,271'b0};
assign c[823913:820896] = {1237'b0,c_w_272,272'b0};
assign c[826931:823914] = {1236'b0,c_w_273,273'b0};
assign c[829949:826932] = {1235'b0,c_w_274,274'b0};
assign c[832967:829950] = {1234'b0,c_w_275,275'b0};
assign c[835985:832968] = {1233'b0,c_w_276,276'b0};
assign c[839003:835986] = {1232'b0,c_w_277,277'b0};
assign c[842021:839004] = {1231'b0,c_w_278,278'b0};
assign c[845039:842022] = {1230'b0,c_w_279,279'b0};
assign c[848057:845040] = {1229'b0,c_w_280,280'b0};
assign c[851075:848058] = {1228'b0,c_w_281,281'b0};
assign c[854093:851076] = {1227'b0,c_w_282,282'b0};
assign c[857111:854094] = {1226'b0,c_w_283,283'b0};
assign c[860129:857112] = {1225'b0,c_w_284,284'b0};
assign c[863147:860130] = {1224'b0,c_w_285,285'b0};
assign c[866165:863148] = {1223'b0,c_w_286,286'b0};
assign c[869183:866166] = {1222'b0,c_w_287,287'b0};
assign c[872201:869184] = {1221'b0,c_w_288,288'b0};
assign c[875219:872202] = {1220'b0,c_w_289,289'b0};
assign c[878237:875220] = {1219'b0,c_w_290,290'b0};
assign c[881255:878238] = {1218'b0,c_w_291,291'b0};
assign c[884273:881256] = {1217'b0,c_w_292,292'b0};
assign c[887291:884274] = {1216'b0,c_w_293,293'b0};
assign c[890309:887292] = {1215'b0,c_w_294,294'b0};
assign c[893327:890310] = {1214'b0,c_w_295,295'b0};
assign c[896345:893328] = {1213'b0,c_w_296,296'b0};
assign c[899363:896346] = {1212'b0,c_w_297,297'b0};
assign c[902381:899364] = {1211'b0,c_w_298,298'b0};
assign c[905399:902382] = {1210'b0,c_w_299,299'b0};
assign c[908417:905400] = {1209'b0,c_w_300,300'b0};
assign c[911435:908418] = {1208'b0,c_w_301,301'b0};
assign c[914453:911436] = {1207'b0,c_w_302,302'b0};
assign c[917471:914454] = {1206'b0,c_w_303,303'b0};
assign c[920489:917472] = {1205'b0,c_w_304,304'b0};
assign c[923507:920490] = {1204'b0,c_w_305,305'b0};
assign c[926525:923508] = {1203'b0,c_w_306,306'b0};
assign c[929543:926526] = {1202'b0,c_w_307,307'b0};
assign c[932561:929544] = {1201'b0,c_w_308,308'b0};
assign c[935579:932562] = {1200'b0,c_w_309,309'b0};
assign c[938597:935580] = {1199'b0,c_w_310,310'b0};
assign c[941615:938598] = {1198'b0,c_w_311,311'b0};
assign c[944633:941616] = {1197'b0,c_w_312,312'b0};
assign c[947651:944634] = {1196'b0,c_w_313,313'b0};
assign c[950669:947652] = {1195'b0,c_w_314,314'b0};
assign c[953687:950670] = {1194'b0,c_w_315,315'b0};
assign c[956705:953688] = {1193'b0,c_w_316,316'b0};
assign c[959723:956706] = {1192'b0,c_w_317,317'b0};
assign c[962741:959724] = {1191'b0,c_w_318,318'b0};
assign c[965759:962742] = {1190'b0,c_w_319,319'b0};
assign c[968777:965760] = {1189'b0,c_w_320,320'b0};
assign c[971795:968778] = {1188'b0,c_w_321,321'b0};
assign c[974813:971796] = {1187'b0,c_w_322,322'b0};
assign c[977831:974814] = {1186'b0,c_w_323,323'b0};
assign c[980849:977832] = {1185'b0,c_w_324,324'b0};
assign c[983867:980850] = {1184'b0,c_w_325,325'b0};
assign c[986885:983868] = {1183'b0,c_w_326,326'b0};
assign c[989903:986886] = {1182'b0,c_w_327,327'b0};
assign c[992921:989904] = {1181'b0,c_w_328,328'b0};
assign c[995939:992922] = {1180'b0,c_w_329,329'b0};
assign c[998957:995940] = {1179'b0,c_w_330,330'b0};
assign c[1001975:998958] = {1178'b0,c_w_331,331'b0};
assign c[1004993:1001976] = {1177'b0,c_w_332,332'b0};
assign c[1008011:1004994] = {1176'b0,c_w_333,333'b0};
assign c[1011029:1008012] = {1175'b0,c_w_334,334'b0};
assign c[1014047:1011030] = {1174'b0,c_w_335,335'b0};
assign c[1017065:1014048] = {1173'b0,c_w_336,336'b0};
assign c[1020083:1017066] = {1172'b0,c_w_337,337'b0};
assign c[1023101:1020084] = {1171'b0,c_w_338,338'b0};
assign c[1026119:1023102] = {1170'b0,c_w_339,339'b0};
assign c[1029137:1026120] = {1169'b0,c_w_340,340'b0};
assign c[1032155:1029138] = {1168'b0,c_w_341,341'b0};
assign c[1035173:1032156] = {1167'b0,c_w_342,342'b0};
assign c[1038191:1035174] = {1166'b0,c_w_343,343'b0};
assign c[1041209:1038192] = {1165'b0,c_w_344,344'b0};
assign c[1044227:1041210] = {1164'b0,c_w_345,345'b0};
assign c[1047245:1044228] = {1163'b0,c_w_346,346'b0};
assign c[1050263:1047246] = {1162'b0,c_w_347,347'b0};
assign c[1053281:1050264] = {1161'b0,c_w_348,348'b0};
assign c[1056299:1053282] = {1160'b0,c_w_349,349'b0};
assign c[1059317:1056300] = {1159'b0,c_w_350,350'b0};
assign c[1062335:1059318] = {1158'b0,c_w_351,351'b0};
assign c[1065353:1062336] = {1157'b0,c_w_352,352'b0};
assign c[1068371:1065354] = {1156'b0,c_w_353,353'b0};
assign c[1071389:1068372] = {1155'b0,c_w_354,354'b0};
assign c[1074407:1071390] = {1154'b0,c_w_355,355'b0};
assign c[1077425:1074408] = {1153'b0,c_w_356,356'b0};
assign c[1080443:1077426] = {1152'b0,c_w_357,357'b0};
assign c[1083461:1080444] = {1151'b0,c_w_358,358'b0};
assign c[1086479:1083462] = {1150'b0,c_w_359,359'b0};
assign c[1089497:1086480] = {1149'b0,c_w_360,360'b0};
assign c[1092515:1089498] = {1148'b0,c_w_361,361'b0};
assign c[1095533:1092516] = {1147'b0,c_w_362,362'b0};
assign c[1098551:1095534] = {1146'b0,c_w_363,363'b0};
assign c[1101569:1098552] = {1145'b0,c_w_364,364'b0};
assign c[1104587:1101570] = {1144'b0,c_w_365,365'b0};
assign c[1107605:1104588] = {1143'b0,c_w_366,366'b0};
assign c[1110623:1107606] = {1142'b0,c_w_367,367'b0};
assign c[1113641:1110624] = {1141'b0,c_w_368,368'b0};
assign c[1116659:1113642] = {1140'b0,c_w_369,369'b0};
assign c[1119677:1116660] = {1139'b0,c_w_370,370'b0};
assign c[1122695:1119678] = {1138'b0,c_w_371,371'b0};
assign c[1125713:1122696] = {1137'b0,c_w_372,372'b0};
assign c[1128731:1125714] = {1136'b0,c_w_373,373'b0};
assign c[1131749:1128732] = {1135'b0,c_w_374,374'b0};
assign c[1134767:1131750] = {1134'b0,c_w_375,375'b0};
assign c[1137785:1134768] = {1133'b0,c_w_376,376'b0};
assign c[1140803:1137786] = {1132'b0,c_w_377,377'b0};
assign c[1143821:1140804] = {1131'b0,c_w_378,378'b0};
assign c[1146839:1143822] = {1130'b0,c_w_379,379'b0};
assign c[1149857:1146840] = {1129'b0,c_w_380,380'b0};
assign c[1152875:1149858] = {1128'b0,c_w_381,381'b0};
assign c[1155893:1152876] = {1127'b0,c_w_382,382'b0};
assign c[1158911:1155894] = {1126'b0,c_w_383,383'b0};
assign c[1161929:1158912] = {1125'b0,c_w_384,384'b0};
assign c[1164947:1161930] = {1124'b0,c_w_385,385'b0};
assign c[1167965:1164948] = {1123'b0,c_w_386,386'b0};
assign c[1170983:1167966] = {1122'b0,c_w_387,387'b0};
assign c[1174001:1170984] = {1121'b0,c_w_388,388'b0};
assign c[1177019:1174002] = {1120'b0,c_w_389,389'b0};
assign c[1180037:1177020] = {1119'b0,c_w_390,390'b0};
assign c[1183055:1180038] = {1118'b0,c_w_391,391'b0};
assign c[1186073:1183056] = {1117'b0,c_w_392,392'b0};
assign c[1189091:1186074] = {1116'b0,c_w_393,393'b0};
assign c[1192109:1189092] = {1115'b0,c_w_394,394'b0};
assign c[1195127:1192110] = {1114'b0,c_w_395,395'b0};
assign c[1198145:1195128] = {1113'b0,c_w_396,396'b0};
assign c[1201163:1198146] = {1112'b0,c_w_397,397'b0};
assign c[1204181:1201164] = {1111'b0,c_w_398,398'b0};
assign c[1207199:1204182] = {1110'b0,c_w_399,399'b0};
assign c[1210217:1207200] = {1109'b0,c_w_400,400'b0};
assign c[1213235:1210218] = {1108'b0,c_w_401,401'b0};
assign c[1216253:1213236] = {1107'b0,c_w_402,402'b0};
assign c[1219271:1216254] = {1106'b0,c_w_403,403'b0};
assign c[1222289:1219272] = {1105'b0,c_w_404,404'b0};
assign c[1225307:1222290] = {1104'b0,c_w_405,405'b0};
assign c[1228325:1225308] = {1103'b0,c_w_406,406'b0};
assign c[1231343:1228326] = {1102'b0,c_w_407,407'b0};
assign c[1234361:1231344] = {1101'b0,c_w_408,408'b0};
assign c[1237379:1234362] = {1100'b0,c_w_409,409'b0};
assign c[1240397:1237380] = {1099'b0,c_w_410,410'b0};
assign c[1243415:1240398] = {1098'b0,c_w_411,411'b0};
assign c[1246433:1243416] = {1097'b0,c_w_412,412'b0};
assign c[1249451:1246434] = {1096'b0,c_w_413,413'b0};
assign c[1252469:1249452] = {1095'b0,c_w_414,414'b0};
assign c[1255487:1252470] = {1094'b0,c_w_415,415'b0};
assign c[1258505:1255488] = {1093'b0,c_w_416,416'b0};
assign c[1261523:1258506] = {1092'b0,c_w_417,417'b0};
assign c[1264541:1261524] = {1091'b0,c_w_418,418'b0};
assign c[1267559:1264542] = {1090'b0,c_w_419,419'b0};
assign c[1270577:1267560] = {1089'b0,c_w_420,420'b0};
assign c[1273595:1270578] = {1088'b0,c_w_421,421'b0};
assign c[1276613:1273596] = {1087'b0,c_w_422,422'b0};
assign c[1279631:1276614] = {1086'b0,c_w_423,423'b0};
assign c[1282649:1279632] = {1085'b0,c_w_424,424'b0};
assign c[1285667:1282650] = {1084'b0,c_w_425,425'b0};
assign c[1288685:1285668] = {1083'b0,c_w_426,426'b0};
assign c[1291703:1288686] = {1082'b0,c_w_427,427'b0};
assign c[1294721:1291704] = {1081'b0,c_w_428,428'b0};
assign c[1297739:1294722] = {1080'b0,c_w_429,429'b0};
assign c[1300757:1297740] = {1079'b0,c_w_430,430'b0};
assign c[1303775:1300758] = {1078'b0,c_w_431,431'b0};
assign c[1306793:1303776] = {1077'b0,c_w_432,432'b0};
assign c[1309811:1306794] = {1076'b0,c_w_433,433'b0};
assign c[1312829:1309812] = {1075'b0,c_w_434,434'b0};
assign c[1315847:1312830] = {1074'b0,c_w_435,435'b0};
assign c[1318865:1315848] = {1073'b0,c_w_436,436'b0};
assign c[1321883:1318866] = {1072'b0,c_w_437,437'b0};
assign c[1324901:1321884] = {1071'b0,c_w_438,438'b0};
assign c[1327919:1324902] = {1070'b0,c_w_439,439'b0};
assign c[1330937:1327920] = {1069'b0,c_w_440,440'b0};
assign c[1333955:1330938] = {1068'b0,c_w_441,441'b0};
assign c[1336973:1333956] = {1067'b0,c_w_442,442'b0};
assign c[1339991:1336974] = {1066'b0,c_w_443,443'b0};
assign c[1343009:1339992] = {1065'b0,c_w_444,444'b0};
assign c[1346027:1343010] = {1064'b0,c_w_445,445'b0};
assign c[1349045:1346028] = {1063'b0,c_w_446,446'b0};
assign c[1352063:1349046] = {1062'b0,c_w_447,447'b0};
assign c[1355081:1352064] = {1061'b0,c_w_448,448'b0};
assign c[1358099:1355082] = {1060'b0,c_w_449,449'b0};
assign c[1361117:1358100] = {1059'b0,c_w_450,450'b0};
assign c[1364135:1361118] = {1058'b0,c_w_451,451'b0};
assign c[1367153:1364136] = {1057'b0,c_w_452,452'b0};
assign c[1370171:1367154] = {1056'b0,c_w_453,453'b0};
assign c[1373189:1370172] = {1055'b0,c_w_454,454'b0};
assign c[1376207:1373190] = {1054'b0,c_w_455,455'b0};
assign c[1379225:1376208] = {1053'b0,c_w_456,456'b0};
assign c[1382243:1379226] = {1052'b0,c_w_457,457'b0};
assign c[1385261:1382244] = {1051'b0,c_w_458,458'b0};
assign c[1388279:1385262] = {1050'b0,c_w_459,459'b0};
assign c[1391297:1388280] = {1049'b0,c_w_460,460'b0};
assign c[1394315:1391298] = {1048'b0,c_w_461,461'b0};
assign c[1397333:1394316] = {1047'b0,c_w_462,462'b0};
assign c[1400351:1397334] = {1046'b0,c_w_463,463'b0};
assign c[1403369:1400352] = {1045'b0,c_w_464,464'b0};
assign c[1406387:1403370] = {1044'b0,c_w_465,465'b0};
assign c[1409405:1406388] = {1043'b0,c_w_466,466'b0};
assign c[1412423:1409406] = {1042'b0,c_w_467,467'b0};
assign c[1415441:1412424] = {1041'b0,c_w_468,468'b0};
assign c[1418459:1415442] = {1040'b0,c_w_469,469'b0};
assign c[1421477:1418460] = {1039'b0,c_w_470,470'b0};
assign c[1424495:1421478] = {1038'b0,c_w_471,471'b0};
assign c[1427513:1424496] = {1037'b0,c_w_472,472'b0};
assign c[1430531:1427514] = {1036'b0,c_w_473,473'b0};
assign c[1433549:1430532] = {1035'b0,c_w_474,474'b0};
assign c[1436567:1433550] = {1034'b0,c_w_475,475'b0};
assign c[1439585:1436568] = {1033'b0,c_w_476,476'b0};
assign c[1442603:1439586] = {1032'b0,c_w_477,477'b0};
assign c[1445621:1442604] = {1031'b0,c_w_478,478'b0};
assign c[1448639:1445622] = {1030'b0,c_w_479,479'b0};
assign c[1451657:1448640] = {1029'b0,c_w_480,480'b0};
assign c[1454675:1451658] = {1028'b0,c_w_481,481'b0};
assign c[1457693:1454676] = {1027'b0,c_w_482,482'b0};
assign c[1460711:1457694] = {1026'b0,c_w_483,483'b0};
assign c[1463729:1460712] = {1025'b0,c_w_484,484'b0};
assign c[1466747:1463730] = {1024'b0,c_w_485,485'b0};
assign c[1469765:1466748] = {1023'b0,c_w_486,486'b0};
assign c[1472783:1469766] = {1022'b0,c_w_487,487'b0};
assign c[1475801:1472784] = {1021'b0,c_w_488,488'b0};
assign c[1478819:1475802] = {1020'b0,c_w_489,489'b0};
assign c[1481837:1478820] = {1019'b0,c_w_490,490'b0};
assign c[1484855:1481838] = {1018'b0,c_w_491,491'b0};
assign c[1487873:1484856] = {1017'b0,c_w_492,492'b0};
assign c[1490891:1487874] = {1016'b0,c_w_493,493'b0};
assign c[1493909:1490892] = {1015'b0,c_w_494,494'b0};
assign c[1496927:1493910] = {1014'b0,c_w_495,495'b0};
assign c[1499945:1496928] = {1013'b0,c_w_496,496'b0};
assign c[1502963:1499946] = {1012'b0,c_w_497,497'b0};
assign c[1505981:1502964] = {1011'b0,c_w_498,498'b0};
assign c[1508999:1505982] = {1010'b0,c_w_499,499'b0};
assign c[1512017:1509000] = {1009'b0,c_w_500,500'b0};
assign c[1515035:1512018] = {1008'b0,c_w_501,501'b0};
assign c[1518053:1515036] = {1007'b0,c_w_502,502'b0};
assign c[1521071:1518054] = {1006'b0,c_w_503,503'b0};
assign c[1524089:1521072] = {1005'b0,c_w_504,504'b0};
assign c[1527107:1524090] = {1004'b0,c_w_505,505'b0};
assign c[1530125:1527108] = {1003'b0,c_w_506,506'b0};
assign c[1533143:1530126] = {1002'b0,c_w_507,507'b0};
assign c[1536161:1533144] = {1001'b0,c_w_508,508'b0};
assign c[1539179:1536162] = {1000'b0,c_w_509,509'b0};
assign c[1542197:1539180] = {999'b0,c_w_510,510'b0};
assign c[1545215:1542198] = {998'b0,c_w_511,511'b0};
assign c[1548233:1545216] = {997'b0,c_w_512,512'b0};
assign c[1551251:1548234] = {996'b0,c_w_513,513'b0};
assign c[1554269:1551252] = {995'b0,c_w_514,514'b0};
assign c[1557287:1554270] = {994'b0,c_w_515,515'b0};
assign c[1560305:1557288] = {993'b0,c_w_516,516'b0};
assign c[1563323:1560306] = {992'b0,c_w_517,517'b0};
assign c[1566341:1563324] = {991'b0,c_w_518,518'b0};
assign c[1569359:1566342] = {990'b0,c_w_519,519'b0};
assign c[1572377:1569360] = {989'b0,c_w_520,520'b0};
assign c[1575395:1572378] = {988'b0,c_w_521,521'b0};
assign c[1578413:1575396] = {987'b0,c_w_522,522'b0};
assign c[1581431:1578414] = {986'b0,c_w_523,523'b0};
assign c[1584449:1581432] = {985'b0,c_w_524,524'b0};
assign c[1587467:1584450] = {984'b0,c_w_525,525'b0};
assign c[1590485:1587468] = {983'b0,c_w_526,526'b0};
assign c[1593503:1590486] = {982'b0,c_w_527,527'b0};
assign c[1596521:1593504] = {981'b0,c_w_528,528'b0};
assign c[1599539:1596522] = {980'b0,c_w_529,529'b0};
assign c[1602557:1599540] = {979'b0,c_w_530,530'b0};
assign c[1605575:1602558] = {978'b0,c_w_531,531'b0};
assign c[1608593:1605576] = {977'b0,c_w_532,532'b0};
assign c[1611611:1608594] = {976'b0,c_w_533,533'b0};
assign c[1614629:1611612] = {975'b0,c_w_534,534'b0};
assign c[1617647:1614630] = {974'b0,c_w_535,535'b0};
assign c[1620665:1617648] = {973'b0,c_w_536,536'b0};
assign c[1623683:1620666] = {972'b0,c_w_537,537'b0};
assign c[1626701:1623684] = {971'b0,c_w_538,538'b0};
assign c[1629719:1626702] = {970'b0,c_w_539,539'b0};
assign c[1632737:1629720] = {969'b0,c_w_540,540'b0};
assign c[1635755:1632738] = {968'b0,c_w_541,541'b0};
assign c[1638773:1635756] = {967'b0,c_w_542,542'b0};
assign c[1641791:1638774] = {966'b0,c_w_543,543'b0};
assign c[1644809:1641792] = {965'b0,c_w_544,544'b0};
assign c[1647827:1644810] = {964'b0,c_w_545,545'b0};
assign c[1650845:1647828] = {963'b0,c_w_546,546'b0};
assign c[1653863:1650846] = {962'b0,c_w_547,547'b0};
assign c[1656881:1653864] = {961'b0,c_w_548,548'b0};
assign c[1659899:1656882] = {960'b0,c_w_549,549'b0};
assign c[1662917:1659900] = {959'b0,c_w_550,550'b0};
assign c[1665935:1662918] = {958'b0,c_w_551,551'b0};
assign c[1668953:1665936] = {957'b0,c_w_552,552'b0};
assign c[1671971:1668954] = {956'b0,c_w_553,553'b0};
assign c[1674989:1671972] = {955'b0,c_w_554,554'b0};
assign c[1678007:1674990] = {954'b0,c_w_555,555'b0};
assign c[1681025:1678008] = {953'b0,c_w_556,556'b0};
assign c[1684043:1681026] = {952'b0,c_w_557,557'b0};
assign c[1687061:1684044] = {951'b0,c_w_558,558'b0};
assign c[1690079:1687062] = {950'b0,c_w_559,559'b0};
assign c[1693097:1690080] = {949'b0,c_w_560,560'b0};
assign c[1696115:1693098] = {948'b0,c_w_561,561'b0};
assign c[1699133:1696116] = {947'b0,c_w_562,562'b0};
assign c[1702151:1699134] = {946'b0,c_w_563,563'b0};
assign c[1705169:1702152] = {945'b0,c_w_564,564'b0};
assign c[1708187:1705170] = {944'b0,c_w_565,565'b0};
assign c[1711205:1708188] = {943'b0,c_w_566,566'b0};
assign c[1714223:1711206] = {942'b0,c_w_567,567'b0};
assign c[1717241:1714224] = {941'b0,c_w_568,568'b0};
assign c[1720259:1717242] = {940'b0,c_w_569,569'b0};
assign c[1723277:1720260] = {939'b0,c_w_570,570'b0};
assign c[1726295:1723278] = {938'b0,c_w_571,571'b0};
assign c[1729313:1726296] = {937'b0,c_w_572,572'b0};
assign c[1732331:1729314] = {936'b0,c_w_573,573'b0};
assign c[1735349:1732332] = {935'b0,c_w_574,574'b0};
assign c[1738367:1735350] = {934'b0,c_w_575,575'b0};
assign c[1741385:1738368] = {933'b0,c_w_576,576'b0};
assign c[1744403:1741386] = {932'b0,c_w_577,577'b0};
assign c[1747421:1744404] = {931'b0,c_w_578,578'b0};
assign c[1750439:1747422] = {930'b0,c_w_579,579'b0};
assign c[1753457:1750440] = {929'b0,c_w_580,580'b0};
assign c[1756475:1753458] = {928'b0,c_w_581,581'b0};
assign c[1759493:1756476] = {927'b0,c_w_582,582'b0};
assign c[1762511:1759494] = {926'b0,c_w_583,583'b0};
assign c[1765529:1762512] = {925'b0,c_w_584,584'b0};
assign c[1768547:1765530] = {924'b0,c_w_585,585'b0};
assign c[1771565:1768548] = {923'b0,c_w_586,586'b0};
assign c[1774583:1771566] = {922'b0,c_w_587,587'b0};
assign c[1777601:1774584] = {921'b0,c_w_588,588'b0};
assign c[1780619:1777602] = {920'b0,c_w_589,589'b0};
assign c[1783637:1780620] = {919'b0,c_w_590,590'b0};
assign c[1786655:1783638] = {918'b0,c_w_591,591'b0};
assign c[1789673:1786656] = {917'b0,c_w_592,592'b0};
assign c[1792691:1789674] = {916'b0,c_w_593,593'b0};
assign c[1795709:1792692] = {915'b0,c_w_594,594'b0};
assign c[1798727:1795710] = {914'b0,c_w_595,595'b0};
assign c[1801745:1798728] = {913'b0,c_w_596,596'b0};
assign c[1804763:1801746] = {912'b0,c_w_597,597'b0};
assign c[1807781:1804764] = {911'b0,c_w_598,598'b0};
assign c[1810799:1807782] = {910'b0,c_w_599,599'b0};
assign c[1813817:1810800] = {909'b0,c_w_600,600'b0};
assign c[1816835:1813818] = {908'b0,c_w_601,601'b0};
assign c[1819853:1816836] = {907'b0,c_w_602,602'b0};
assign c[1822871:1819854] = {906'b0,c_w_603,603'b0};
assign c[1825889:1822872] = {905'b0,c_w_604,604'b0};
assign c[1828907:1825890] = {904'b0,c_w_605,605'b0};
assign c[1831925:1828908] = {903'b0,c_w_606,606'b0};
assign c[1834943:1831926] = {902'b0,c_w_607,607'b0};
assign c[1837961:1834944] = {901'b0,c_w_608,608'b0};
assign c[1840979:1837962] = {900'b0,c_w_609,609'b0};
assign c[1843997:1840980] = {899'b0,c_w_610,610'b0};
assign c[1847015:1843998] = {898'b0,c_w_611,611'b0};
assign c[1850033:1847016] = {897'b0,c_w_612,612'b0};
assign c[1853051:1850034] = {896'b0,c_w_613,613'b0};
assign c[1856069:1853052] = {895'b0,c_w_614,614'b0};
assign c[1859087:1856070] = {894'b0,c_w_615,615'b0};
assign c[1862105:1859088] = {893'b0,c_w_616,616'b0};
assign c[1865123:1862106] = {892'b0,c_w_617,617'b0};
assign c[1868141:1865124] = {891'b0,c_w_618,618'b0};
assign c[1871159:1868142] = {890'b0,c_w_619,619'b0};
assign c[1874177:1871160] = {889'b0,c_w_620,620'b0};
assign c[1877195:1874178] = {888'b0,c_w_621,621'b0};
assign c[1880213:1877196] = {887'b0,c_w_622,622'b0};
assign c[1883231:1880214] = {886'b0,c_w_623,623'b0};
assign c[1886249:1883232] = {885'b0,c_w_624,624'b0};
assign c[1889267:1886250] = {884'b0,c_w_625,625'b0};
assign c[1892285:1889268] = {883'b0,c_w_626,626'b0};
assign c[1895303:1892286] = {882'b0,c_w_627,627'b0};
assign c[1898321:1895304] = {881'b0,c_w_628,628'b0};
assign c[1901339:1898322] = {880'b0,c_w_629,629'b0};
assign c[1904357:1901340] = {879'b0,c_w_630,630'b0};
assign c[1907375:1904358] = {878'b0,c_w_631,631'b0};
assign c[1910393:1907376] = {877'b0,c_w_632,632'b0};
assign c[1913411:1910394] = {876'b0,c_w_633,633'b0};
assign c[1916429:1913412] = {875'b0,c_w_634,634'b0};
assign c[1919447:1916430] = {874'b0,c_w_635,635'b0};
assign c[1922465:1919448] = {873'b0,c_w_636,636'b0};
assign c[1925483:1922466] = {872'b0,c_w_637,637'b0};
assign c[1928501:1925484] = {871'b0,c_w_638,638'b0};
assign c[1931519:1928502] = {870'b0,c_w_639,639'b0};
assign c[1934537:1931520] = {869'b0,c_w_640,640'b0};
assign c[1937555:1934538] = {868'b0,c_w_641,641'b0};
assign c[1940573:1937556] = {867'b0,c_w_642,642'b0};
assign c[1943591:1940574] = {866'b0,c_w_643,643'b0};
assign c[1946609:1943592] = {865'b0,c_w_644,644'b0};
assign c[1949627:1946610] = {864'b0,c_w_645,645'b0};
assign c[1952645:1949628] = {863'b0,c_w_646,646'b0};
assign c[1955663:1952646] = {862'b0,c_w_647,647'b0};
assign c[1958681:1955664] = {861'b0,c_w_648,648'b0};
assign c[1961699:1958682] = {860'b0,c_w_649,649'b0};
assign c[1964717:1961700] = {859'b0,c_w_650,650'b0};
assign c[1967735:1964718] = {858'b0,c_w_651,651'b0};
assign c[1970753:1967736] = {857'b0,c_w_652,652'b0};
assign c[1973771:1970754] = {856'b0,c_w_653,653'b0};
assign c[1976789:1973772] = {855'b0,c_w_654,654'b0};
assign c[1979807:1976790] = {854'b0,c_w_655,655'b0};
assign c[1982825:1979808] = {853'b0,c_w_656,656'b0};
assign c[1985843:1982826] = {852'b0,c_w_657,657'b0};
assign c[1988861:1985844] = {851'b0,c_w_658,658'b0};
assign c[1991879:1988862] = {850'b0,c_w_659,659'b0};
assign c[1994897:1991880] = {849'b0,c_w_660,660'b0};
assign c[1997915:1994898] = {848'b0,c_w_661,661'b0};
assign c[2000933:1997916] = {847'b0,c_w_662,662'b0};
assign c[2003951:2000934] = {846'b0,c_w_663,663'b0};
assign c[2006969:2003952] = {845'b0,c_w_664,664'b0};
assign c[2009987:2006970] = {844'b0,c_w_665,665'b0};
assign c[2013005:2009988] = {843'b0,c_w_666,666'b0};
assign c[2016023:2013006] = {842'b0,c_w_667,667'b0};
assign c[2019041:2016024] = {841'b0,c_w_668,668'b0};
assign c[2022059:2019042] = {840'b0,c_w_669,669'b0};
assign c[2025077:2022060] = {839'b0,c_w_670,670'b0};
assign c[2028095:2025078] = {838'b0,c_w_671,671'b0};
assign c[2031113:2028096] = {837'b0,c_w_672,672'b0};
assign c[2034131:2031114] = {836'b0,c_w_673,673'b0};
assign c[2037149:2034132] = {835'b0,c_w_674,674'b0};
assign c[2040167:2037150] = {834'b0,c_w_675,675'b0};
assign c[2043185:2040168] = {833'b0,c_w_676,676'b0};
assign c[2046203:2043186] = {832'b0,c_w_677,677'b0};
assign c[2049221:2046204] = {831'b0,c_w_678,678'b0};
assign c[2052239:2049222] = {830'b0,c_w_679,679'b0};
assign c[2055257:2052240] = {829'b0,c_w_680,680'b0};
assign c[2058275:2055258] = {828'b0,c_w_681,681'b0};
assign c[2061293:2058276] = {827'b0,c_w_682,682'b0};
assign c[2064311:2061294] = {826'b0,c_w_683,683'b0};
assign c[2067329:2064312] = {825'b0,c_w_684,684'b0};
assign c[2070347:2067330] = {824'b0,c_w_685,685'b0};
assign c[2073365:2070348] = {823'b0,c_w_686,686'b0};
assign c[2076383:2073366] = {822'b0,c_w_687,687'b0};
assign c[2079401:2076384] = {821'b0,c_w_688,688'b0};
assign c[2082419:2079402] = {820'b0,c_w_689,689'b0};
assign c[2085437:2082420] = {819'b0,c_w_690,690'b0};
assign c[2088455:2085438] = {818'b0,c_w_691,691'b0};
assign c[2091473:2088456] = {817'b0,c_w_692,692'b0};
assign c[2094491:2091474] = {816'b0,c_w_693,693'b0};
assign c[2097509:2094492] = {815'b0,c_w_694,694'b0};
assign c[2100527:2097510] = {814'b0,c_w_695,695'b0};
assign c[2103545:2100528] = {813'b0,c_w_696,696'b0};
assign c[2106563:2103546] = {812'b0,c_w_697,697'b0};
assign c[2109581:2106564] = {811'b0,c_w_698,698'b0};
assign c[2112599:2109582] = {810'b0,c_w_699,699'b0};
assign c[2115617:2112600] = {809'b0,c_w_700,700'b0};
assign c[2118635:2115618] = {808'b0,c_w_701,701'b0};
assign c[2121653:2118636] = {807'b0,c_w_702,702'b0};
assign c[2124671:2121654] = {806'b0,c_w_703,703'b0};
assign c[2127689:2124672] = {805'b0,c_w_704,704'b0};
assign c[2130707:2127690] = {804'b0,c_w_705,705'b0};
assign c[2133725:2130708] = {803'b0,c_w_706,706'b0};
assign c[2136743:2133726] = {802'b0,c_w_707,707'b0};
assign c[2139761:2136744] = {801'b0,c_w_708,708'b0};
assign c[2142779:2139762] = {800'b0,c_w_709,709'b0};
assign c[2145797:2142780] = {799'b0,c_w_710,710'b0};
assign c[2148815:2145798] = {798'b0,c_w_711,711'b0};
assign c[2151833:2148816] = {797'b0,c_w_712,712'b0};
assign c[2154851:2151834] = {796'b0,c_w_713,713'b0};
assign c[2157869:2154852] = {795'b0,c_w_714,714'b0};
assign c[2160887:2157870] = {794'b0,c_w_715,715'b0};
assign c[2163905:2160888] = {793'b0,c_w_716,716'b0};
assign c[2166923:2163906] = {792'b0,c_w_717,717'b0};
assign c[2169941:2166924] = {791'b0,c_w_718,718'b0};
assign c[2172959:2169942] = {790'b0,c_w_719,719'b0};
assign c[2175977:2172960] = {789'b0,c_w_720,720'b0};
assign c[2178995:2175978] = {788'b0,c_w_721,721'b0};
assign c[2182013:2178996] = {787'b0,c_w_722,722'b0};
assign c[2185031:2182014] = {786'b0,c_w_723,723'b0};
assign c[2188049:2185032] = {785'b0,c_w_724,724'b0};
assign c[2191067:2188050] = {784'b0,c_w_725,725'b0};
assign c[2194085:2191068] = {783'b0,c_w_726,726'b0};
assign c[2197103:2194086] = {782'b0,c_w_727,727'b0};
assign c[2200121:2197104] = {781'b0,c_w_728,728'b0};
assign c[2203139:2200122] = {780'b0,c_w_729,729'b0};
assign c[2206157:2203140] = {779'b0,c_w_730,730'b0};
assign c[2209175:2206158] = {778'b0,c_w_731,731'b0};
assign c[2212193:2209176] = {777'b0,c_w_732,732'b0};
assign c[2215211:2212194] = {776'b0,c_w_733,733'b0};
assign c[2218229:2215212] = {775'b0,c_w_734,734'b0};
assign c[2221247:2218230] = {774'b0,c_w_735,735'b0};
assign c[2224265:2221248] = {773'b0,c_w_736,736'b0};
assign c[2227283:2224266] = {772'b0,c_w_737,737'b0};
assign c[2230301:2227284] = {771'b0,c_w_738,738'b0};
assign c[2233319:2230302] = {770'b0,c_w_739,739'b0};
assign c[2236337:2233320] = {769'b0,c_w_740,740'b0};
assign c[2239355:2236338] = {768'b0,c_w_741,741'b0};
assign c[2242373:2239356] = {767'b0,c_w_742,742'b0};
assign c[2245391:2242374] = {766'b0,c_w_743,743'b0};
assign c[2248409:2245392] = {765'b0,c_w_744,744'b0};
assign c[2251427:2248410] = {764'b0,c_w_745,745'b0};
assign c[2254445:2251428] = {763'b0,c_w_746,746'b0};
assign c[2257463:2254446] = {762'b0,c_w_747,747'b0};
assign c[2260481:2257464] = {761'b0,c_w_748,748'b0};
assign c[2263499:2260482] = {760'b0,c_w_749,749'b0};
assign c[2266517:2263500] = {759'b0,c_w_750,750'b0};
assign c[2269535:2266518] = {758'b0,c_w_751,751'b0};
assign c[2272553:2269536] = {757'b0,c_w_752,752'b0};
assign c[2275571:2272554] = {756'b0,c_w_753,753'b0};
assign c[2278589:2275572] = {755'b0,c_w_754,754'b0};
assign c[2281607:2278590] = {754'b0,c_w_755,755'b0};
assign c[2284625:2281608] = {753'b0,c_w_756,756'b0};
assign c[2287643:2284626] = {752'b0,c_w_757,757'b0};
assign c[2290661:2287644] = {751'b0,c_w_758,758'b0};
assign c[2293679:2290662] = {750'b0,c_w_759,759'b0};
assign c[2296697:2293680] = {749'b0,c_w_760,760'b0};
assign c[2299715:2296698] = {748'b0,c_w_761,761'b0};
assign c[2302733:2299716] = {747'b0,c_w_762,762'b0};
assign c[2305751:2302734] = {746'b0,c_w_763,763'b0};
assign c[2308769:2305752] = {745'b0,c_w_764,764'b0};
assign c[2311787:2308770] = {744'b0,c_w_765,765'b0};
assign c[2314805:2311788] = {743'b0,c_w_766,766'b0};
assign c[2317823:2314806] = {742'b0,c_w_767,767'b0};
assign c[2320841:2317824] = {741'b0,c_w_768,768'b0};
assign c[2323859:2320842] = {740'b0,c_w_769,769'b0};
assign c[2326877:2323860] = {739'b0,c_w_770,770'b0};
assign c[2329895:2326878] = {738'b0,c_w_771,771'b0};
assign c[2332913:2329896] = {737'b0,c_w_772,772'b0};
assign c[2335931:2332914] = {736'b0,c_w_773,773'b0};
assign c[2338949:2335932] = {735'b0,c_w_774,774'b0};
assign c[2341967:2338950] = {734'b0,c_w_775,775'b0};
assign c[2344985:2341968] = {733'b0,c_w_776,776'b0};
assign c[2348003:2344986] = {732'b0,c_w_777,777'b0};
assign c[2351021:2348004] = {731'b0,c_w_778,778'b0};
assign c[2354039:2351022] = {730'b0,c_w_779,779'b0};
assign c[2357057:2354040] = {729'b0,c_w_780,780'b0};
assign c[2360075:2357058] = {728'b0,c_w_781,781'b0};
assign c[2363093:2360076] = {727'b0,c_w_782,782'b0};
assign c[2366111:2363094] = {726'b0,c_w_783,783'b0};
assign c[2369129:2366112] = {725'b0,c_w_784,784'b0};
assign c[2372147:2369130] = {724'b0,c_w_785,785'b0};
assign c[2375165:2372148] = {723'b0,c_w_786,786'b0};
assign c[2378183:2375166] = {722'b0,c_w_787,787'b0};
assign c[2381201:2378184] = {721'b0,c_w_788,788'b0};
assign c[2384219:2381202] = {720'b0,c_w_789,789'b0};
assign c[2387237:2384220] = {719'b0,c_w_790,790'b0};
assign c[2390255:2387238] = {718'b0,c_w_791,791'b0};
assign c[2393273:2390256] = {717'b0,c_w_792,792'b0};
assign c[2396291:2393274] = {716'b0,c_w_793,793'b0};
assign c[2399309:2396292] = {715'b0,c_w_794,794'b0};
assign c[2402327:2399310] = {714'b0,c_w_795,795'b0};
assign c[2405345:2402328] = {713'b0,c_w_796,796'b0};
assign c[2408363:2405346] = {712'b0,c_w_797,797'b0};
assign c[2411381:2408364] = {711'b0,c_w_798,798'b0};
assign c[2414399:2411382] = {710'b0,c_w_799,799'b0};
assign c[2417417:2414400] = {709'b0,c_w_800,800'b0};
assign c[2420435:2417418] = {708'b0,c_w_801,801'b0};
assign c[2423453:2420436] = {707'b0,c_w_802,802'b0};
assign c[2426471:2423454] = {706'b0,c_w_803,803'b0};
assign c[2429489:2426472] = {705'b0,c_w_804,804'b0};
assign c[2432507:2429490] = {704'b0,c_w_805,805'b0};
assign c[2435525:2432508] = {703'b0,c_w_806,806'b0};
assign c[2438543:2435526] = {702'b0,c_w_807,807'b0};
assign c[2441561:2438544] = {701'b0,c_w_808,808'b0};
assign c[2444579:2441562] = {700'b0,c_w_809,809'b0};
assign c[2447597:2444580] = {699'b0,c_w_810,810'b0};
assign c[2450615:2447598] = {698'b0,c_w_811,811'b0};
assign c[2453633:2450616] = {697'b0,c_w_812,812'b0};
assign c[2456651:2453634] = {696'b0,c_w_813,813'b0};
assign c[2459669:2456652] = {695'b0,c_w_814,814'b0};
assign c[2462687:2459670] = {694'b0,c_w_815,815'b0};
assign c[2465705:2462688] = {693'b0,c_w_816,816'b0};
assign c[2468723:2465706] = {692'b0,c_w_817,817'b0};
assign c[2471741:2468724] = {691'b0,c_w_818,818'b0};
assign c[2474759:2471742] = {690'b0,c_w_819,819'b0};
assign c[2477777:2474760] = {689'b0,c_w_820,820'b0};
assign c[2480795:2477778] = {688'b0,c_w_821,821'b0};
assign c[2483813:2480796] = {687'b0,c_w_822,822'b0};
assign c[2486831:2483814] = {686'b0,c_w_823,823'b0};
assign c[2489849:2486832] = {685'b0,c_w_824,824'b0};
assign c[2492867:2489850] = {684'b0,c_w_825,825'b0};
assign c[2495885:2492868] = {683'b0,c_w_826,826'b0};
assign c[2498903:2495886] = {682'b0,c_w_827,827'b0};
assign c[2501921:2498904] = {681'b0,c_w_828,828'b0};
assign c[2504939:2501922] = {680'b0,c_w_829,829'b0};
assign c[2507957:2504940] = {679'b0,c_w_830,830'b0};
assign c[2510975:2507958] = {678'b0,c_w_831,831'b0};
assign c[2513993:2510976] = {677'b0,c_w_832,832'b0};
assign c[2517011:2513994] = {676'b0,c_w_833,833'b0};
assign c[2520029:2517012] = {675'b0,c_w_834,834'b0};
assign c[2523047:2520030] = {674'b0,c_w_835,835'b0};
assign c[2526065:2523048] = {673'b0,c_w_836,836'b0};
assign c[2529083:2526066] = {672'b0,c_w_837,837'b0};
assign c[2532101:2529084] = {671'b0,c_w_838,838'b0};
assign c[2535119:2532102] = {670'b0,c_w_839,839'b0};
assign c[2538137:2535120] = {669'b0,c_w_840,840'b0};
assign c[2541155:2538138] = {668'b0,c_w_841,841'b0};
assign c[2544173:2541156] = {667'b0,c_w_842,842'b0};
assign c[2547191:2544174] = {666'b0,c_w_843,843'b0};
assign c[2550209:2547192] = {665'b0,c_w_844,844'b0};
assign c[2553227:2550210] = {664'b0,c_w_845,845'b0};
assign c[2556245:2553228] = {663'b0,c_w_846,846'b0};
assign c[2559263:2556246] = {662'b0,c_w_847,847'b0};
assign c[2562281:2559264] = {661'b0,c_w_848,848'b0};
assign c[2565299:2562282] = {660'b0,c_w_849,849'b0};
assign c[2568317:2565300] = {659'b0,c_w_850,850'b0};
assign c[2571335:2568318] = {658'b0,c_w_851,851'b0};
assign c[2574353:2571336] = {657'b0,c_w_852,852'b0};
assign c[2577371:2574354] = {656'b0,c_w_853,853'b0};
assign c[2580389:2577372] = {655'b0,c_w_854,854'b0};
assign c[2583407:2580390] = {654'b0,c_w_855,855'b0};
assign c[2586425:2583408] = {653'b0,c_w_856,856'b0};
assign c[2589443:2586426] = {652'b0,c_w_857,857'b0};
assign c[2592461:2589444] = {651'b0,c_w_858,858'b0};
assign c[2595479:2592462] = {650'b0,c_w_859,859'b0};
assign c[2598497:2595480] = {649'b0,c_w_860,860'b0};
assign c[2601515:2598498] = {648'b0,c_w_861,861'b0};
assign c[2604533:2601516] = {647'b0,c_w_862,862'b0};
assign c[2607551:2604534] = {646'b0,c_w_863,863'b0};
assign c[2610569:2607552] = {645'b0,c_w_864,864'b0};
assign c[2613587:2610570] = {644'b0,c_w_865,865'b0};
assign c[2616605:2613588] = {643'b0,c_w_866,866'b0};
assign c[2619623:2616606] = {642'b0,c_w_867,867'b0};
assign c[2622641:2619624] = {641'b0,c_w_868,868'b0};
assign c[2625659:2622642] = {640'b0,c_w_869,869'b0};
assign c[2628677:2625660] = {639'b0,c_w_870,870'b0};
assign c[2631695:2628678] = {638'b0,c_w_871,871'b0};
assign c[2634713:2631696] = {637'b0,c_w_872,872'b0};
assign c[2637731:2634714] = {636'b0,c_w_873,873'b0};
assign c[2640749:2637732] = {635'b0,c_w_874,874'b0};
assign c[2643767:2640750] = {634'b0,c_w_875,875'b0};
assign c[2646785:2643768] = {633'b0,c_w_876,876'b0};
assign c[2649803:2646786] = {632'b0,c_w_877,877'b0};
assign c[2652821:2649804] = {631'b0,c_w_878,878'b0};
assign c[2655839:2652822] = {630'b0,c_w_879,879'b0};
assign c[2658857:2655840] = {629'b0,c_w_880,880'b0};
assign c[2661875:2658858] = {628'b0,c_w_881,881'b0};
assign c[2664893:2661876] = {627'b0,c_w_882,882'b0};
assign c[2667911:2664894] = {626'b0,c_w_883,883'b0};
assign c[2670929:2667912] = {625'b0,c_w_884,884'b0};
assign c[2673947:2670930] = {624'b0,c_w_885,885'b0};
assign c[2676965:2673948] = {623'b0,c_w_886,886'b0};
assign c[2679983:2676966] = {622'b0,c_w_887,887'b0};
assign c[2683001:2679984] = {621'b0,c_w_888,888'b0};
assign c[2686019:2683002] = {620'b0,c_w_889,889'b0};
assign c[2689037:2686020] = {619'b0,c_w_890,890'b0};
assign c[2692055:2689038] = {618'b0,c_w_891,891'b0};
assign c[2695073:2692056] = {617'b0,c_w_892,892'b0};
assign c[2698091:2695074] = {616'b0,c_w_893,893'b0};
assign c[2701109:2698092] = {615'b0,c_w_894,894'b0};
assign c[2704127:2701110] = {614'b0,c_w_895,895'b0};
assign c[2707145:2704128] = {613'b0,c_w_896,896'b0};
assign c[2710163:2707146] = {612'b0,c_w_897,897'b0};
assign c[2713181:2710164] = {611'b0,c_w_898,898'b0};
assign c[2716199:2713182] = {610'b0,c_w_899,899'b0};
assign c[2719217:2716200] = {609'b0,c_w_900,900'b0};
assign c[2722235:2719218] = {608'b0,c_w_901,901'b0};
assign c[2725253:2722236] = {607'b0,c_w_902,902'b0};
assign c[2728271:2725254] = {606'b0,c_w_903,903'b0};
assign c[2731289:2728272] = {605'b0,c_w_904,904'b0};
assign c[2734307:2731290] = {604'b0,c_w_905,905'b0};
assign c[2737325:2734308] = {603'b0,c_w_906,906'b0};
assign c[2740343:2737326] = {602'b0,c_w_907,907'b0};
assign c[2743361:2740344] = {601'b0,c_w_908,908'b0};
assign c[2746379:2743362] = {600'b0,c_w_909,909'b0};
assign c[2749397:2746380] = {599'b0,c_w_910,910'b0};
assign c[2752415:2749398] = {598'b0,c_w_911,911'b0};
assign c[2755433:2752416] = {597'b0,c_w_912,912'b0};
assign c[2758451:2755434] = {596'b0,c_w_913,913'b0};
assign c[2761469:2758452] = {595'b0,c_w_914,914'b0};
assign c[2764487:2761470] = {594'b0,c_w_915,915'b0};
assign c[2767505:2764488] = {593'b0,c_w_916,916'b0};
assign c[2770523:2767506] = {592'b0,c_w_917,917'b0};
assign c[2773541:2770524] = {591'b0,c_w_918,918'b0};
assign c[2776559:2773542] = {590'b0,c_w_919,919'b0};
assign c[2779577:2776560] = {589'b0,c_w_920,920'b0};
assign c[2782595:2779578] = {588'b0,c_w_921,921'b0};
assign c[2785613:2782596] = {587'b0,c_w_922,922'b0};
assign c[2788631:2785614] = {586'b0,c_w_923,923'b0};
assign c[2791649:2788632] = {585'b0,c_w_924,924'b0};
assign c[2794667:2791650] = {584'b0,c_w_925,925'b0};
assign c[2797685:2794668] = {583'b0,c_w_926,926'b0};
assign c[2800703:2797686] = {582'b0,c_w_927,927'b0};
assign c[2803721:2800704] = {581'b0,c_w_928,928'b0};
assign c[2806739:2803722] = {580'b0,c_w_929,929'b0};
assign c[2809757:2806740] = {579'b0,c_w_930,930'b0};
assign c[2812775:2809758] = {578'b0,c_w_931,931'b0};
assign c[2815793:2812776] = {577'b0,c_w_932,932'b0};
assign c[2818811:2815794] = {576'b0,c_w_933,933'b0};
assign c[2821829:2818812] = {575'b0,c_w_934,934'b0};
assign c[2824847:2821830] = {574'b0,c_w_935,935'b0};
assign c[2827865:2824848] = {573'b0,c_w_936,936'b0};
assign c[2830883:2827866] = {572'b0,c_w_937,937'b0};
assign c[2833901:2830884] = {571'b0,c_w_938,938'b0};
assign c[2836919:2833902] = {570'b0,c_w_939,939'b0};
assign c[2839937:2836920] = {569'b0,c_w_940,940'b0};
assign c[2842955:2839938] = {568'b0,c_w_941,941'b0};
assign c[2845973:2842956] = {567'b0,c_w_942,942'b0};
assign c[2848991:2845974] = {566'b0,c_w_943,943'b0};
assign c[2852009:2848992] = {565'b0,c_w_944,944'b0};
assign c[2855027:2852010] = {564'b0,c_w_945,945'b0};
assign c[2858045:2855028] = {563'b0,c_w_946,946'b0};
assign c[2861063:2858046] = {562'b0,c_w_947,947'b0};
assign c[2864081:2861064] = {561'b0,c_w_948,948'b0};
assign c[2867099:2864082] = {560'b0,c_w_949,949'b0};
assign c[2870117:2867100] = {559'b0,c_w_950,950'b0};
assign c[2873135:2870118] = {558'b0,c_w_951,951'b0};
assign c[2876153:2873136] = {557'b0,c_w_952,952'b0};
assign c[2879171:2876154] = {556'b0,c_w_953,953'b0};
assign c[2882189:2879172] = {555'b0,c_w_954,954'b0};
assign c[2885207:2882190] = {554'b0,c_w_955,955'b0};
assign c[2888225:2885208] = {553'b0,c_w_956,956'b0};
assign c[2891243:2888226] = {552'b0,c_w_957,957'b0};
assign c[2894261:2891244] = {551'b0,c_w_958,958'b0};
assign c[2897279:2894262] = {550'b0,c_w_959,959'b0};
assign c[2900297:2897280] = {549'b0,c_w_960,960'b0};
assign c[2903315:2900298] = {548'b0,c_w_961,961'b0};
assign c[2906333:2903316] = {547'b0,c_w_962,962'b0};
assign c[2909351:2906334] = {546'b0,c_w_963,963'b0};
assign c[2912369:2909352] = {545'b0,c_w_964,964'b0};
assign c[2915387:2912370] = {544'b0,c_w_965,965'b0};
assign c[2918405:2915388] = {543'b0,c_w_966,966'b0};
assign c[2921423:2918406] = {542'b0,c_w_967,967'b0};
assign c[2924441:2921424] = {541'b0,c_w_968,968'b0};
assign c[2927459:2924442] = {540'b0,c_w_969,969'b0};
assign c[2930477:2927460] = {539'b0,c_w_970,970'b0};
assign c[2933495:2930478] = {538'b0,c_w_971,971'b0};
assign c[2936513:2933496] = {537'b0,c_w_972,972'b0};
assign c[2939531:2936514] = {536'b0,c_w_973,973'b0};
assign c[2942549:2939532] = {535'b0,c_w_974,974'b0};
assign c[2945567:2942550] = {534'b0,c_w_975,975'b0};
assign c[2948585:2945568] = {533'b0,c_w_976,976'b0};
assign c[2951603:2948586] = {532'b0,c_w_977,977'b0};
assign c[2954621:2951604] = {531'b0,c_w_978,978'b0};
assign c[2957639:2954622] = {530'b0,c_w_979,979'b0};
assign c[2960657:2957640] = {529'b0,c_w_980,980'b0};
assign c[2963675:2960658] = {528'b0,c_w_981,981'b0};
assign c[2966693:2963676] = {527'b0,c_w_982,982'b0};
assign c[2969711:2966694] = {526'b0,c_w_983,983'b0};
assign c[2972729:2969712] = {525'b0,c_w_984,984'b0};
assign c[2975747:2972730] = {524'b0,c_w_985,985'b0};
assign c[2978765:2975748] = {523'b0,c_w_986,986'b0};
assign c[2981783:2978766] = {522'b0,c_w_987,987'b0};
assign c[2984801:2981784] = {521'b0,c_w_988,988'b0};
assign c[2987819:2984802] = {520'b0,c_w_989,989'b0};
assign c[2990837:2987820] = {519'b0,c_w_990,990'b0};
assign c[2993855:2990838] = {518'b0,c_w_991,991'b0};
assign c[2996873:2993856] = {517'b0,c_w_992,992'b0};
assign c[2999891:2996874] = {516'b0,c_w_993,993'b0};
assign c[3002909:2999892] = {515'b0,c_w_994,994'b0};
assign c[3005927:3002910] = {514'b0,c_w_995,995'b0};
assign c[3008945:3005928] = {513'b0,c_w_996,996'b0};
assign c[3011963:3008946] = {512'b0,c_w_997,997'b0};
assign c[3014981:3011964] = {511'b0,c_w_998,998'b0};
assign c[3017999:3014982] = {510'b0,c_w_999,999'b0};
assign c[3021017:3018000] = {509'b0,c_w_1000,1000'b0};
assign c[3024035:3021018] = {508'b0,c_w_1001,1001'b0};
assign c[3027053:3024036] = {507'b0,c_w_1002,1002'b0};
assign c[3030071:3027054] = {506'b0,c_w_1003,1003'b0};
assign c[3033089:3030072] = {505'b0,c_w_1004,1004'b0};
assign c[3036107:3033090] = {504'b0,c_w_1005,1005'b0};
assign c[3039125:3036108] = {503'b0,c_w_1006,1006'b0};
assign c[3042143:3039126] = {502'b0,c_w_1007,1007'b0};
assign c[3045161:3042144] = {501'b0,c_w_1008,1008'b0};
assign c[3048179:3045162] = {500'b0,c_w_1009,1009'b0};
assign c[3051197:3048180] = {499'b0,c_w_1010,1010'b0};
assign c[3054215:3051198] = {498'b0,c_w_1011,1011'b0};
assign c[3057233:3054216] = {497'b0,c_w_1012,1012'b0};
assign c[3060251:3057234] = {496'b0,c_w_1013,1013'b0};
assign c[3063269:3060252] = {495'b0,c_w_1014,1014'b0};
assign c[3066287:3063270] = {494'b0,c_w_1015,1015'b0};
assign c[3069305:3066288] = {493'b0,c_w_1016,1016'b0};
assign c[3072323:3069306] = {492'b0,c_w_1017,1017'b0};
assign c[3075341:3072324] = {491'b0,c_w_1018,1018'b0};
assign c[3078359:3075342] = {490'b0,c_w_1019,1019'b0};
assign c[3081377:3078360] = {489'b0,c_w_1020,1020'b0};
assign c[3084395:3081378] = {488'b0,c_w_1021,1021'b0};
assign c[3087413:3084396] = {487'b0,c_w_1022,1022'b0};
assign c[3090431:3087414] = {486'b0,c_w_1023,1023'b0};
assign c[3093449:3090432] = {485'b0,c_w_1024,1024'b0};
assign c[3096467:3093450] = {484'b0,c_w_1025,1025'b0};
assign c[3099485:3096468] = {483'b0,c_w_1026,1026'b0};
assign c[3102503:3099486] = {482'b0,c_w_1027,1027'b0};
assign c[3105521:3102504] = {481'b0,c_w_1028,1028'b0};
assign c[3108539:3105522] = {480'b0,c_w_1029,1029'b0};
assign c[3111557:3108540] = {479'b0,c_w_1030,1030'b0};
assign c[3114575:3111558] = {478'b0,c_w_1031,1031'b0};
assign c[3117593:3114576] = {477'b0,c_w_1032,1032'b0};
assign c[3120611:3117594] = {476'b0,c_w_1033,1033'b0};
assign c[3123629:3120612] = {475'b0,c_w_1034,1034'b0};
assign c[3126647:3123630] = {474'b0,c_w_1035,1035'b0};
assign c[3129665:3126648] = {473'b0,c_w_1036,1036'b0};
assign c[3132683:3129666] = {472'b0,c_w_1037,1037'b0};
assign c[3135701:3132684] = {471'b0,c_w_1038,1038'b0};
assign c[3138719:3135702] = {470'b0,c_w_1039,1039'b0};
assign c[3141737:3138720] = {469'b0,c_w_1040,1040'b0};
assign c[3144755:3141738] = {468'b0,c_w_1041,1041'b0};
assign c[3147773:3144756] = {467'b0,c_w_1042,1042'b0};
assign c[3150791:3147774] = {466'b0,c_w_1043,1043'b0};
assign c[3153809:3150792] = {465'b0,c_w_1044,1044'b0};
assign c[3156827:3153810] = {464'b0,c_w_1045,1045'b0};
assign c[3159845:3156828] = {463'b0,c_w_1046,1046'b0};
assign c[3162863:3159846] = {462'b0,c_w_1047,1047'b0};
assign c[3165881:3162864] = {461'b0,c_w_1048,1048'b0};
assign c[3168899:3165882] = {460'b0,c_w_1049,1049'b0};
assign c[3171917:3168900] = {459'b0,c_w_1050,1050'b0};
assign c[3174935:3171918] = {458'b0,c_w_1051,1051'b0};
assign c[3177953:3174936] = {457'b0,c_w_1052,1052'b0};
assign c[3180971:3177954] = {456'b0,c_w_1053,1053'b0};
assign c[3183989:3180972] = {455'b0,c_w_1054,1054'b0};
assign c[3187007:3183990] = {454'b0,c_w_1055,1055'b0};
assign c[3190025:3187008] = {453'b0,c_w_1056,1056'b0};
assign c[3193043:3190026] = {452'b0,c_w_1057,1057'b0};
assign c[3196061:3193044] = {451'b0,c_w_1058,1058'b0};
assign c[3199079:3196062] = {450'b0,c_w_1059,1059'b0};
assign c[3202097:3199080] = {449'b0,c_w_1060,1060'b0};
assign c[3205115:3202098] = {448'b0,c_w_1061,1061'b0};
assign c[3208133:3205116] = {447'b0,c_w_1062,1062'b0};
assign c[3211151:3208134] = {446'b0,c_w_1063,1063'b0};
assign c[3214169:3211152] = {445'b0,c_w_1064,1064'b0};
assign c[3217187:3214170] = {444'b0,c_w_1065,1065'b0};
assign c[3220205:3217188] = {443'b0,c_w_1066,1066'b0};
assign c[3223223:3220206] = {442'b0,c_w_1067,1067'b0};
assign c[3226241:3223224] = {441'b0,c_w_1068,1068'b0};
assign c[3229259:3226242] = {440'b0,c_w_1069,1069'b0};
assign c[3232277:3229260] = {439'b0,c_w_1070,1070'b0};
assign c[3235295:3232278] = {438'b0,c_w_1071,1071'b0};
assign c[3238313:3235296] = {437'b0,c_w_1072,1072'b0};
assign c[3241331:3238314] = {436'b0,c_w_1073,1073'b0};
assign c[3244349:3241332] = {435'b0,c_w_1074,1074'b0};
assign c[3247367:3244350] = {434'b0,c_w_1075,1075'b0};
assign c[3250385:3247368] = {433'b0,c_w_1076,1076'b0};
assign c[3253403:3250386] = {432'b0,c_w_1077,1077'b0};
assign c[3256421:3253404] = {431'b0,c_w_1078,1078'b0};
assign c[3259439:3256422] = {430'b0,c_w_1079,1079'b0};
assign c[3262457:3259440] = {429'b0,c_w_1080,1080'b0};
assign c[3265475:3262458] = {428'b0,c_w_1081,1081'b0};
assign c[3268493:3265476] = {427'b0,c_w_1082,1082'b0};
assign c[3271511:3268494] = {426'b0,c_w_1083,1083'b0};
assign c[3274529:3271512] = {425'b0,c_w_1084,1084'b0};
assign c[3277547:3274530] = {424'b0,c_w_1085,1085'b0};
assign c[3280565:3277548] = {423'b0,c_w_1086,1086'b0};
assign c[3283583:3280566] = {422'b0,c_w_1087,1087'b0};
assign c[3286601:3283584] = {421'b0,c_w_1088,1088'b0};
assign c[3289619:3286602] = {420'b0,c_w_1089,1089'b0};
assign c[3292637:3289620] = {419'b0,c_w_1090,1090'b0};
assign c[3295655:3292638] = {418'b0,c_w_1091,1091'b0};
assign c[3298673:3295656] = {417'b0,c_w_1092,1092'b0};
assign c[3301691:3298674] = {416'b0,c_w_1093,1093'b0};
assign c[3304709:3301692] = {415'b0,c_w_1094,1094'b0};
assign c[3307727:3304710] = {414'b0,c_w_1095,1095'b0};
assign c[3310745:3307728] = {413'b0,c_w_1096,1096'b0};
assign c[3313763:3310746] = {412'b0,c_w_1097,1097'b0};
assign c[3316781:3313764] = {411'b0,c_w_1098,1098'b0};
assign c[3319799:3316782] = {410'b0,c_w_1099,1099'b0};
assign c[3322817:3319800] = {409'b0,c_w_1100,1100'b0};
assign c[3325835:3322818] = {408'b0,c_w_1101,1101'b0};
assign c[3328853:3325836] = {407'b0,c_w_1102,1102'b0};
assign c[3331871:3328854] = {406'b0,c_w_1103,1103'b0};
assign c[3334889:3331872] = {405'b0,c_w_1104,1104'b0};
assign c[3337907:3334890] = {404'b0,c_w_1105,1105'b0};
assign c[3340925:3337908] = {403'b0,c_w_1106,1106'b0};
assign c[3343943:3340926] = {402'b0,c_w_1107,1107'b0};
assign c[3346961:3343944] = {401'b0,c_w_1108,1108'b0};
assign c[3349979:3346962] = {400'b0,c_w_1109,1109'b0};
assign c[3352997:3349980] = {399'b0,c_w_1110,1110'b0};
assign c[3356015:3352998] = {398'b0,c_w_1111,1111'b0};
assign c[3359033:3356016] = {397'b0,c_w_1112,1112'b0};
assign c[3362051:3359034] = {396'b0,c_w_1113,1113'b0};
assign c[3365069:3362052] = {395'b0,c_w_1114,1114'b0};
assign c[3368087:3365070] = {394'b0,c_w_1115,1115'b0};
assign c[3371105:3368088] = {393'b0,c_w_1116,1116'b0};
assign c[3374123:3371106] = {392'b0,c_w_1117,1117'b0};
assign c[3377141:3374124] = {391'b0,c_w_1118,1118'b0};
assign c[3380159:3377142] = {390'b0,c_w_1119,1119'b0};
assign c[3383177:3380160] = {389'b0,c_w_1120,1120'b0};
assign c[3386195:3383178] = {388'b0,c_w_1121,1121'b0};
assign c[3389213:3386196] = {387'b0,c_w_1122,1122'b0};
assign c[3392231:3389214] = {386'b0,c_w_1123,1123'b0};
assign c[3395249:3392232] = {385'b0,c_w_1124,1124'b0};
assign c[3398267:3395250] = {384'b0,c_w_1125,1125'b0};
assign c[3401285:3398268] = {383'b0,c_w_1126,1126'b0};
assign c[3404303:3401286] = {382'b0,c_w_1127,1127'b0};
assign c[3407321:3404304] = {381'b0,c_w_1128,1128'b0};
assign c[3410339:3407322] = {380'b0,c_w_1129,1129'b0};
assign c[3413357:3410340] = {379'b0,c_w_1130,1130'b0};
assign c[3416375:3413358] = {378'b0,c_w_1131,1131'b0};
assign c[3419393:3416376] = {377'b0,c_w_1132,1132'b0};
assign c[3422411:3419394] = {376'b0,c_w_1133,1133'b0};
assign c[3425429:3422412] = {375'b0,c_w_1134,1134'b0};
assign c[3428447:3425430] = {374'b0,c_w_1135,1135'b0};
assign c[3431465:3428448] = {373'b0,c_w_1136,1136'b0};
assign c[3434483:3431466] = {372'b0,c_w_1137,1137'b0};
assign c[3437501:3434484] = {371'b0,c_w_1138,1138'b0};
assign c[3440519:3437502] = {370'b0,c_w_1139,1139'b0};
assign c[3443537:3440520] = {369'b0,c_w_1140,1140'b0};
assign c[3446555:3443538] = {368'b0,c_w_1141,1141'b0};
assign c[3449573:3446556] = {367'b0,c_w_1142,1142'b0};
assign c[3452591:3449574] = {366'b0,c_w_1143,1143'b0};
assign c[3455609:3452592] = {365'b0,c_w_1144,1144'b0};
assign c[3458627:3455610] = {364'b0,c_w_1145,1145'b0};
assign c[3461645:3458628] = {363'b0,c_w_1146,1146'b0};
assign c[3464663:3461646] = {362'b0,c_w_1147,1147'b0};
assign c[3467681:3464664] = {361'b0,c_w_1148,1148'b0};
assign c[3470699:3467682] = {360'b0,c_w_1149,1149'b0};
assign c[3473717:3470700] = {359'b0,c_w_1150,1150'b0};
assign c[3476735:3473718] = {358'b0,c_w_1151,1151'b0};
assign c[3479753:3476736] = {357'b0,c_w_1152,1152'b0};
assign c[3482771:3479754] = {356'b0,c_w_1153,1153'b0};
assign c[3485789:3482772] = {355'b0,c_w_1154,1154'b0};
assign c[3488807:3485790] = {354'b0,c_w_1155,1155'b0};
assign c[3491825:3488808] = {353'b0,c_w_1156,1156'b0};
assign c[3494843:3491826] = {352'b0,c_w_1157,1157'b0};
assign c[3497861:3494844] = {351'b0,c_w_1158,1158'b0};
assign c[3500879:3497862] = {350'b0,c_w_1159,1159'b0};
assign c[3503897:3500880] = {349'b0,c_w_1160,1160'b0};
assign c[3506915:3503898] = {348'b0,c_w_1161,1161'b0};
assign c[3509933:3506916] = {347'b0,c_w_1162,1162'b0};
assign c[3512951:3509934] = {346'b0,c_w_1163,1163'b0};
assign c[3515969:3512952] = {345'b0,c_w_1164,1164'b0};
assign c[3518987:3515970] = {344'b0,c_w_1165,1165'b0};
assign c[3522005:3518988] = {343'b0,c_w_1166,1166'b0};
assign c[3525023:3522006] = {342'b0,c_w_1167,1167'b0};
assign c[3528041:3525024] = {341'b0,c_w_1168,1168'b0};
assign c[3531059:3528042] = {340'b0,c_w_1169,1169'b0};
assign c[3534077:3531060] = {339'b0,c_w_1170,1170'b0};
assign c[3537095:3534078] = {338'b0,c_w_1171,1171'b0};
assign c[3540113:3537096] = {337'b0,c_w_1172,1172'b0};
assign c[3543131:3540114] = {336'b0,c_w_1173,1173'b0};
assign c[3546149:3543132] = {335'b0,c_w_1174,1174'b0};
assign c[3549167:3546150] = {334'b0,c_w_1175,1175'b0};
assign c[3552185:3549168] = {333'b0,c_w_1176,1176'b0};
assign c[3555203:3552186] = {332'b0,c_w_1177,1177'b0};
assign c[3558221:3555204] = {331'b0,c_w_1178,1178'b0};
assign c[3561239:3558222] = {330'b0,c_w_1179,1179'b0};
assign c[3564257:3561240] = {329'b0,c_w_1180,1180'b0};
assign c[3567275:3564258] = {328'b0,c_w_1181,1181'b0};
assign c[3570293:3567276] = {327'b0,c_w_1182,1182'b0};
assign c[3573311:3570294] = {326'b0,c_w_1183,1183'b0};
assign c[3576329:3573312] = {325'b0,c_w_1184,1184'b0};
assign c[3579347:3576330] = {324'b0,c_w_1185,1185'b0};
assign c[3582365:3579348] = {323'b0,c_w_1186,1186'b0};
assign c[3585383:3582366] = {322'b0,c_w_1187,1187'b0};
assign c[3588401:3585384] = {321'b0,c_w_1188,1188'b0};
assign c[3591419:3588402] = {320'b0,c_w_1189,1189'b0};
assign c[3594437:3591420] = {319'b0,c_w_1190,1190'b0};
assign c[3597455:3594438] = {318'b0,c_w_1191,1191'b0};
assign c[3600473:3597456] = {317'b0,c_w_1192,1192'b0};
assign c[3603491:3600474] = {316'b0,c_w_1193,1193'b0};
assign c[3606509:3603492] = {315'b0,c_w_1194,1194'b0};
assign c[3609527:3606510] = {314'b0,c_w_1195,1195'b0};
assign c[3612545:3609528] = {313'b0,c_w_1196,1196'b0};
assign c[3615563:3612546] = {312'b0,c_w_1197,1197'b0};
assign c[3618581:3615564] = {311'b0,c_w_1198,1198'b0};
assign c[3621599:3618582] = {310'b0,c_w_1199,1199'b0};
assign c[3624617:3621600] = {309'b0,c_w_1200,1200'b0};
assign c[3627635:3624618] = {308'b0,c_w_1201,1201'b0};
assign c[3630653:3627636] = {307'b0,c_w_1202,1202'b0};
assign c[3633671:3630654] = {306'b0,c_w_1203,1203'b0};
assign c[3636689:3633672] = {305'b0,c_w_1204,1204'b0};
assign c[3639707:3636690] = {304'b0,c_w_1205,1205'b0};
assign c[3642725:3639708] = {303'b0,c_w_1206,1206'b0};
assign c[3645743:3642726] = {302'b0,c_w_1207,1207'b0};
assign c[3648761:3645744] = {301'b0,c_w_1208,1208'b0};
assign c[3651779:3648762] = {300'b0,c_w_1209,1209'b0};
assign c[3654797:3651780] = {299'b0,c_w_1210,1210'b0};
assign c[3657815:3654798] = {298'b0,c_w_1211,1211'b0};
assign c[3660833:3657816] = {297'b0,c_w_1212,1212'b0};
assign c[3663851:3660834] = {296'b0,c_w_1213,1213'b0};
assign c[3666869:3663852] = {295'b0,c_w_1214,1214'b0};
assign c[3669887:3666870] = {294'b0,c_w_1215,1215'b0};
assign c[3672905:3669888] = {293'b0,c_w_1216,1216'b0};
assign c[3675923:3672906] = {292'b0,c_w_1217,1217'b0};
assign c[3678941:3675924] = {291'b0,c_w_1218,1218'b0};
assign c[3681959:3678942] = {290'b0,c_w_1219,1219'b0};
assign c[3684977:3681960] = {289'b0,c_w_1220,1220'b0};
assign c[3687995:3684978] = {288'b0,c_w_1221,1221'b0};
assign c[3691013:3687996] = {287'b0,c_w_1222,1222'b0};
assign c[3694031:3691014] = {286'b0,c_w_1223,1223'b0};
assign c[3697049:3694032] = {285'b0,c_w_1224,1224'b0};
assign c[3700067:3697050] = {284'b0,c_w_1225,1225'b0};
assign c[3703085:3700068] = {283'b0,c_w_1226,1226'b0};
assign c[3706103:3703086] = {282'b0,c_w_1227,1227'b0};
assign c[3709121:3706104] = {281'b0,c_w_1228,1228'b0};
assign c[3712139:3709122] = {280'b0,c_w_1229,1229'b0};
assign c[3715157:3712140] = {279'b0,c_w_1230,1230'b0};
assign c[3718175:3715158] = {278'b0,c_w_1231,1231'b0};
assign c[3721193:3718176] = {277'b0,c_w_1232,1232'b0};
assign c[3724211:3721194] = {276'b0,c_w_1233,1233'b0};
assign c[3727229:3724212] = {275'b0,c_w_1234,1234'b0};
assign c[3730247:3727230] = {274'b0,c_w_1235,1235'b0};
assign c[3733265:3730248] = {273'b0,c_w_1236,1236'b0};
assign c[3736283:3733266] = {272'b0,c_w_1237,1237'b0};
assign c[3739301:3736284] = {271'b0,c_w_1238,1238'b0};
assign c[3742319:3739302] = {270'b0,c_w_1239,1239'b0};
assign c[3745337:3742320] = {269'b0,c_w_1240,1240'b0};
assign c[3748355:3745338] = {268'b0,c_w_1241,1241'b0};
assign c[3751373:3748356] = {267'b0,c_w_1242,1242'b0};
assign c[3754391:3751374] = {266'b0,c_w_1243,1243'b0};
assign c[3757409:3754392] = {265'b0,c_w_1244,1244'b0};
assign c[3760427:3757410] = {264'b0,c_w_1245,1245'b0};
assign c[3763445:3760428] = {263'b0,c_w_1246,1246'b0};
assign c[3766463:3763446] = {262'b0,c_w_1247,1247'b0};
assign c[3769481:3766464] = {261'b0,c_w_1248,1248'b0};
assign c[3772499:3769482] = {260'b0,c_w_1249,1249'b0};
assign c[3775517:3772500] = {259'b0,c_w_1250,1250'b0};
assign c[3778535:3775518] = {258'b0,c_w_1251,1251'b0};
assign c[3781553:3778536] = {257'b0,c_w_1252,1252'b0};
assign c[3784571:3781554] = {256'b0,c_w_1253,1253'b0};
assign c[3787589:3784572] = {255'b0,c_w_1254,1254'b0};
assign c[3790607:3787590] = {254'b0,c_w_1255,1255'b0};
assign c[3793625:3790608] = {253'b0,c_w_1256,1256'b0};
assign c[3796643:3793626] = {252'b0,c_w_1257,1257'b0};
assign c[3799661:3796644] = {251'b0,c_w_1258,1258'b0};
assign c[3802679:3799662] = {250'b0,c_w_1259,1259'b0};
assign c[3805697:3802680] = {249'b0,c_w_1260,1260'b0};
assign c[3808715:3805698] = {248'b0,c_w_1261,1261'b0};
assign c[3811733:3808716] = {247'b0,c_w_1262,1262'b0};
assign c[3814751:3811734] = {246'b0,c_w_1263,1263'b0};
assign c[3817769:3814752] = {245'b0,c_w_1264,1264'b0};
assign c[3820787:3817770] = {244'b0,c_w_1265,1265'b0};
assign c[3823805:3820788] = {243'b0,c_w_1266,1266'b0};
assign c[3826823:3823806] = {242'b0,c_w_1267,1267'b0};
assign c[3829841:3826824] = {241'b0,c_w_1268,1268'b0};
assign c[3832859:3829842] = {240'b0,c_w_1269,1269'b0};
assign c[3835877:3832860] = {239'b0,c_w_1270,1270'b0};
assign c[3838895:3835878] = {238'b0,c_w_1271,1271'b0};
assign c[3841913:3838896] = {237'b0,c_w_1272,1272'b0};
assign c[3844931:3841914] = {236'b0,c_w_1273,1273'b0};
assign c[3847949:3844932] = {235'b0,c_w_1274,1274'b0};
assign c[3850967:3847950] = {234'b0,c_w_1275,1275'b0};
assign c[3853985:3850968] = {233'b0,c_w_1276,1276'b0};
assign c[3857003:3853986] = {232'b0,c_w_1277,1277'b0};
assign c[3860021:3857004] = {231'b0,c_w_1278,1278'b0};
assign c[3863039:3860022] = {230'b0,c_w_1279,1279'b0};
assign c[3866057:3863040] = {229'b0,c_w_1280,1280'b0};
assign c[3869075:3866058] = {228'b0,c_w_1281,1281'b0};
assign c[3872093:3869076] = {227'b0,c_w_1282,1282'b0};
assign c[3875111:3872094] = {226'b0,c_w_1283,1283'b0};
assign c[3878129:3875112] = {225'b0,c_w_1284,1284'b0};
assign c[3881147:3878130] = {224'b0,c_w_1285,1285'b0};
assign c[3884165:3881148] = {223'b0,c_w_1286,1286'b0};
assign c[3887183:3884166] = {222'b0,c_w_1287,1287'b0};
assign c[3890201:3887184] = {221'b0,c_w_1288,1288'b0};
assign c[3893219:3890202] = {220'b0,c_w_1289,1289'b0};
assign c[3896237:3893220] = {219'b0,c_w_1290,1290'b0};
assign c[3899255:3896238] = {218'b0,c_w_1291,1291'b0};
assign c[3902273:3899256] = {217'b0,c_w_1292,1292'b0};
assign c[3905291:3902274] = {216'b0,c_w_1293,1293'b0};
assign c[3908309:3905292] = {215'b0,c_w_1294,1294'b0};
assign c[3911327:3908310] = {214'b0,c_w_1295,1295'b0};
assign c[3914345:3911328] = {213'b0,c_w_1296,1296'b0};
assign c[3917363:3914346] = {212'b0,c_w_1297,1297'b0};
assign c[3920381:3917364] = {211'b0,c_w_1298,1298'b0};
assign c[3923399:3920382] = {210'b0,c_w_1299,1299'b0};
assign c[3926417:3923400] = {209'b0,c_w_1300,1300'b0};
assign c[3929435:3926418] = {208'b0,c_w_1301,1301'b0};
assign c[3932453:3929436] = {207'b0,c_w_1302,1302'b0};
assign c[3935471:3932454] = {206'b0,c_w_1303,1303'b0};
assign c[3938489:3935472] = {205'b0,c_w_1304,1304'b0};
assign c[3941507:3938490] = {204'b0,c_w_1305,1305'b0};
assign c[3944525:3941508] = {203'b0,c_w_1306,1306'b0};
assign c[3947543:3944526] = {202'b0,c_w_1307,1307'b0};
assign c[3950561:3947544] = {201'b0,c_w_1308,1308'b0};
assign c[3953579:3950562] = {200'b0,c_w_1309,1309'b0};
assign c[3956597:3953580] = {199'b0,c_w_1310,1310'b0};
assign c[3959615:3956598] = {198'b0,c_w_1311,1311'b0};
assign c[3962633:3959616] = {197'b0,c_w_1312,1312'b0};
assign c[3965651:3962634] = {196'b0,c_w_1313,1313'b0};
assign c[3968669:3965652] = {195'b0,c_w_1314,1314'b0};
assign c[3971687:3968670] = {194'b0,c_w_1315,1315'b0};
assign c[3974705:3971688] = {193'b0,c_w_1316,1316'b0};
assign c[3977723:3974706] = {192'b0,c_w_1317,1317'b0};
assign c[3980741:3977724] = {191'b0,c_w_1318,1318'b0};
assign c[3983759:3980742] = {190'b0,c_w_1319,1319'b0};
assign c[3986777:3983760] = {189'b0,c_w_1320,1320'b0};
assign c[3989795:3986778] = {188'b0,c_w_1321,1321'b0};
assign c[3992813:3989796] = {187'b0,c_w_1322,1322'b0};
assign c[3995831:3992814] = {186'b0,c_w_1323,1323'b0};
assign c[3998849:3995832] = {185'b0,c_w_1324,1324'b0};
assign c[4001867:3998850] = {184'b0,c_w_1325,1325'b0};
assign c[4004885:4001868] = {183'b0,c_w_1326,1326'b0};
assign c[4007903:4004886] = {182'b0,c_w_1327,1327'b0};
assign c[4010921:4007904] = {181'b0,c_w_1328,1328'b0};
assign c[4013939:4010922] = {180'b0,c_w_1329,1329'b0};
assign c[4016957:4013940] = {179'b0,c_w_1330,1330'b0};
assign c[4019975:4016958] = {178'b0,c_w_1331,1331'b0};
assign c[4022993:4019976] = {177'b0,c_w_1332,1332'b0};
assign c[4026011:4022994] = {176'b0,c_w_1333,1333'b0};
assign c[4029029:4026012] = {175'b0,c_w_1334,1334'b0};
assign c[4032047:4029030] = {174'b0,c_w_1335,1335'b0};
assign c[4035065:4032048] = {173'b0,c_w_1336,1336'b0};
assign c[4038083:4035066] = {172'b0,c_w_1337,1337'b0};
assign c[4041101:4038084] = {171'b0,c_w_1338,1338'b0};
assign c[4044119:4041102] = {170'b0,c_w_1339,1339'b0};
assign c[4047137:4044120] = {169'b0,c_w_1340,1340'b0};
assign c[4050155:4047138] = {168'b0,c_w_1341,1341'b0};
assign c[4053173:4050156] = {167'b0,c_w_1342,1342'b0};
assign c[4056191:4053174] = {166'b0,c_w_1343,1343'b0};
assign c[4059209:4056192] = {165'b0,c_w_1344,1344'b0};
assign c[4062227:4059210] = {164'b0,c_w_1345,1345'b0};
assign c[4065245:4062228] = {163'b0,c_w_1346,1346'b0};
assign c[4068263:4065246] = {162'b0,c_w_1347,1347'b0};
assign c[4071281:4068264] = {161'b0,c_w_1348,1348'b0};
assign c[4074299:4071282] = {160'b0,c_w_1349,1349'b0};
assign c[4077317:4074300] = {159'b0,c_w_1350,1350'b0};
assign c[4080335:4077318] = {158'b0,c_w_1351,1351'b0};
assign c[4083353:4080336] = {157'b0,c_w_1352,1352'b0};
assign c[4086371:4083354] = {156'b0,c_w_1353,1353'b0};
assign c[4089389:4086372] = {155'b0,c_w_1354,1354'b0};
assign c[4092407:4089390] = {154'b0,c_w_1355,1355'b0};
assign c[4095425:4092408] = {153'b0,c_w_1356,1356'b0};
assign c[4098443:4095426] = {152'b0,c_w_1357,1357'b0};
assign c[4101461:4098444] = {151'b0,c_w_1358,1358'b0};
assign c[4104479:4101462] = {150'b0,c_w_1359,1359'b0};
assign c[4107497:4104480] = {149'b0,c_w_1360,1360'b0};
assign c[4110515:4107498] = {148'b0,c_w_1361,1361'b0};
assign c[4113533:4110516] = {147'b0,c_w_1362,1362'b0};
assign c[4116551:4113534] = {146'b0,c_w_1363,1363'b0};
assign c[4119569:4116552] = {145'b0,c_w_1364,1364'b0};
assign c[4122587:4119570] = {144'b0,c_w_1365,1365'b0};
assign c[4125605:4122588] = {143'b0,c_w_1366,1366'b0};
assign c[4128623:4125606] = {142'b0,c_w_1367,1367'b0};
assign c[4131641:4128624] = {141'b0,c_w_1368,1368'b0};
assign c[4134659:4131642] = {140'b0,c_w_1369,1369'b0};
assign c[4137677:4134660] = {139'b0,c_w_1370,1370'b0};
assign c[4140695:4137678] = {138'b0,c_w_1371,1371'b0};
assign c[4143713:4140696] = {137'b0,c_w_1372,1372'b0};
assign c[4146731:4143714] = {136'b0,c_w_1373,1373'b0};
assign c[4149749:4146732] = {135'b0,c_w_1374,1374'b0};
assign c[4152767:4149750] = {134'b0,c_w_1375,1375'b0};
assign c[4155785:4152768] = {133'b0,c_w_1376,1376'b0};
assign c[4158803:4155786] = {132'b0,c_w_1377,1377'b0};
assign c[4161821:4158804] = {131'b0,c_w_1378,1378'b0};
assign c[4164839:4161822] = {130'b0,c_w_1379,1379'b0};
assign c[4167857:4164840] = {129'b0,c_w_1380,1380'b0};
assign c[4170875:4167858] = {128'b0,c_w_1381,1381'b0};
assign c[4173893:4170876] = {127'b0,c_w_1382,1382'b0};
assign c[4176911:4173894] = {126'b0,c_w_1383,1383'b0};
assign c[4179929:4176912] = {125'b0,c_w_1384,1384'b0};
assign c[4182947:4179930] = {124'b0,c_w_1385,1385'b0};
assign c[4185965:4182948] = {123'b0,c_w_1386,1386'b0};
assign c[4188983:4185966] = {122'b0,c_w_1387,1387'b0};
assign c[4192001:4188984] = {121'b0,c_w_1388,1388'b0};
assign c[4195019:4192002] = {120'b0,c_w_1389,1389'b0};
assign c[4198037:4195020] = {119'b0,c_w_1390,1390'b0};
assign c[4201055:4198038] = {118'b0,c_w_1391,1391'b0};
assign c[4204073:4201056] = {117'b0,c_w_1392,1392'b0};
assign c[4207091:4204074] = {116'b0,c_w_1393,1393'b0};
assign c[4210109:4207092] = {115'b0,c_w_1394,1394'b0};
assign c[4213127:4210110] = {114'b0,c_w_1395,1395'b0};
assign c[4216145:4213128] = {113'b0,c_w_1396,1396'b0};
assign c[4219163:4216146] = {112'b0,c_w_1397,1397'b0};
assign c[4222181:4219164] = {111'b0,c_w_1398,1398'b0};
assign c[4225199:4222182] = {110'b0,c_w_1399,1399'b0};
assign c[4228217:4225200] = {109'b0,c_w_1400,1400'b0};
assign c[4231235:4228218] = {108'b0,c_w_1401,1401'b0};
assign c[4234253:4231236] = {107'b0,c_w_1402,1402'b0};
assign c[4237271:4234254] = {106'b0,c_w_1403,1403'b0};
assign c[4240289:4237272] = {105'b0,c_w_1404,1404'b0};
assign c[4243307:4240290] = {104'b0,c_w_1405,1405'b0};
assign c[4246325:4243308] = {103'b0,c_w_1406,1406'b0};
assign c[4249343:4246326] = {102'b0,c_w_1407,1407'b0};
assign c[4252361:4249344] = {101'b0,c_w_1408,1408'b0};
assign c[4255379:4252362] = {100'b0,c_w_1409,1409'b0};
assign c[4258397:4255380] = {99'b0,c_w_1410,1410'b0};
assign c[4261415:4258398] = {98'b0,c_w_1411,1411'b0};
assign c[4264433:4261416] = {97'b0,c_w_1412,1412'b0};
assign c[4267451:4264434] = {96'b0,c_w_1413,1413'b0};
assign c[4270469:4267452] = {95'b0,c_w_1414,1414'b0};
assign c[4273487:4270470] = {94'b0,c_w_1415,1415'b0};
assign c[4276505:4273488] = {93'b0,c_w_1416,1416'b0};
assign c[4279523:4276506] = {92'b0,c_w_1417,1417'b0};
assign c[4282541:4279524] = {91'b0,c_w_1418,1418'b0};
assign c[4285559:4282542] = {90'b0,c_w_1419,1419'b0};
assign c[4288577:4285560] = {89'b0,c_w_1420,1420'b0};
assign c[4291595:4288578] = {88'b0,c_w_1421,1421'b0};
assign c[4294613:4291596] = {87'b0,c_w_1422,1422'b0};
assign c[4297631:4294614] = {86'b0,c_w_1423,1423'b0};
assign c[4300649:4297632] = {85'b0,c_w_1424,1424'b0};
assign c[4303667:4300650] = {84'b0,c_w_1425,1425'b0};
assign c[4306685:4303668] = {83'b0,c_w_1426,1426'b0};
assign c[4309703:4306686] = {82'b0,c_w_1427,1427'b0};
assign c[4312721:4309704] = {81'b0,c_w_1428,1428'b0};
assign c[4315739:4312722] = {80'b0,c_w_1429,1429'b0};
assign c[4318757:4315740] = {79'b0,c_w_1430,1430'b0};
assign c[4321775:4318758] = {78'b0,c_w_1431,1431'b0};
assign c[4324793:4321776] = {77'b0,c_w_1432,1432'b0};
assign c[4327811:4324794] = {76'b0,c_w_1433,1433'b0};
assign c[4330829:4327812] = {75'b0,c_w_1434,1434'b0};
assign c[4333847:4330830] = {74'b0,c_w_1435,1435'b0};
assign c[4336865:4333848] = {73'b0,c_w_1436,1436'b0};
assign c[4339883:4336866] = {72'b0,c_w_1437,1437'b0};
assign c[4342901:4339884] = {71'b0,c_w_1438,1438'b0};
assign c[4345919:4342902] = {70'b0,c_w_1439,1439'b0};
assign c[4348937:4345920] = {69'b0,c_w_1440,1440'b0};
assign c[4351955:4348938] = {68'b0,c_w_1441,1441'b0};
assign c[4354973:4351956] = {67'b0,c_w_1442,1442'b0};
assign c[4357991:4354974] = {66'b0,c_w_1443,1443'b0};
assign c[4361009:4357992] = {65'b0,c_w_1444,1444'b0};
assign c[4364027:4361010] = {64'b0,c_w_1445,1445'b0};
assign c[4367045:4364028] = {63'b0,c_w_1446,1446'b0};
assign c[4370063:4367046] = {62'b0,c_w_1447,1447'b0};
assign c[4373081:4370064] = {61'b0,c_w_1448,1448'b0};
assign c[4376099:4373082] = {60'b0,c_w_1449,1449'b0};
assign c[4379117:4376100] = {59'b0,c_w_1450,1450'b0};
assign c[4382135:4379118] = {58'b0,c_w_1451,1451'b0};
assign c[4385153:4382136] = {57'b0,c_w_1452,1452'b0};
assign c[4388171:4385154] = {56'b0,c_w_1453,1453'b0};
assign c[4391189:4388172] = {55'b0,c_w_1454,1454'b0};
assign c[4394207:4391190] = {54'b0,c_w_1455,1455'b0};
assign c[4397225:4394208] = {53'b0,c_w_1456,1456'b0};
assign c[4400243:4397226] = {52'b0,c_w_1457,1457'b0};
assign c[4403261:4400244] = {51'b0,c_w_1458,1458'b0};
assign c[4406279:4403262] = {50'b0,c_w_1459,1459'b0};
assign c[4409297:4406280] = {49'b0,c_w_1460,1460'b0};
assign c[4412315:4409298] = {48'b0,c_w_1461,1461'b0};
assign c[4415333:4412316] = {47'b0,c_w_1462,1462'b0};
assign c[4418351:4415334] = {46'b0,c_w_1463,1463'b0};
assign c[4421369:4418352] = {45'b0,c_w_1464,1464'b0};
assign c[4424387:4421370] = {44'b0,c_w_1465,1465'b0};
assign c[4427405:4424388] = {43'b0,c_w_1466,1466'b0};
assign c[4430423:4427406] = {42'b0,c_w_1467,1467'b0};
assign c[4433441:4430424] = {41'b0,c_w_1468,1468'b0};
assign c[4436459:4433442] = {40'b0,c_w_1469,1469'b0};
assign c[4439477:4436460] = {39'b0,c_w_1470,1470'b0};
assign c[4442495:4439478] = {38'b0,c_w_1471,1471'b0};
assign c[4445513:4442496] = {37'b0,c_w_1472,1472'b0};
assign c[4448531:4445514] = {36'b0,c_w_1473,1473'b0};
assign c[4451549:4448532] = {35'b0,c_w_1474,1474'b0};
assign c[4454567:4451550] = {34'b0,c_w_1475,1475'b0};
assign c[4457585:4454568] = {33'b0,c_w_1476,1476'b0};
assign c[4460603:4457586] = {32'b0,c_w_1477,1477'b0};
assign c[4463621:4460604] = {31'b0,c_w_1478,1478'b0};
assign c[4466639:4463622] = {30'b0,c_w_1479,1479'b0};
assign c[4469657:4466640] = {29'b0,c_w_1480,1480'b0};
assign c[4472675:4469658] = {28'b0,c_w_1481,1481'b0};
assign c[4475693:4472676] = {27'b0,c_w_1482,1482'b0};
assign c[4478711:4475694] = {26'b0,c_w_1483,1483'b0};
assign c[4481729:4478712] = {25'b0,c_w_1484,1484'b0};
assign c[4484747:4481730] = {24'b0,c_w_1485,1485'b0};
assign c[4487765:4484748] = {23'b0,c_w_1486,1486'b0};
assign c[4490783:4487766] = {22'b0,c_w_1487,1487'b0};
assign c[4493801:4490784] = {21'b0,c_w_1488,1488'b0};
assign c[4496819:4493802] = {20'b0,c_w_1489,1489'b0};
assign c[4499837:4496820] = {19'b0,c_w_1490,1490'b0};
assign c[4502855:4499838] = {18'b0,c_w_1491,1491'b0};
assign c[4505873:4502856] = {17'b0,c_w_1492,1492'b0};
assign c[4508891:4505874] = {16'b0,c_w_1493,1493'b0};
assign c[4511909:4508892] = {15'b0,c_w_1494,1494'b0};
assign c[4514927:4511910] = {14'b0,c_w_1495,1495'b0};
assign c[4517945:4514928] = {13'b0,c_w_1496,1496'b0};
assign c[4520963:4517946] = {12'b0,c_w_1497,1497'b0};
assign c[4523981:4520964] = {11'b0,c_w_1498,1498'b0};
assign c[4526999:4523982] = {10'b0,c_w_1499,1499'b0};
assign c[4530017:4527000] = {9'b0,c_w_1500,1500'b0};
assign c[4533035:4530018] = {8'b0,c_w_1501,1501'b0};
assign c[4536053:4533036] = {7'b0,c_w_1502,1502'b0};
assign c[4539071:4536054] = {6'b0,c_w_1503,1503'b0};
assign c[4542089:4539072] = {5'b0,c_w_1504,1504'b0};
assign c[4545107:4542090] = {4'b0,c_w_1505,1505'b0};
assign c[4548125:4545108] = {3'b0,c_w_1506,1506'b0};
assign c[4551143:4548126] = {2'b0,c_w_1507,1507'b0};
assign c[4554161:4551144] = {1'b0,c_w_1508,1508'b0};
    
endmodule
    